##
## LEF for PtnCells ;
## created by Innovus v19.12-s087_1 on Fri Dec 20 18:37:05 2024
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MLP_no_sram
  CLASS BLOCK ;
  SIZE 368.980000 BY 437.570000 ;
  FOREIGN MLP_no_sram 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 5.065000 0.000000 5.205000 0.140000 ;
    END
  END clk
  PIN rst_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 6.745000 0.000000 6.885000 0.140000 ;
    END
  END rst_b
  PIN start_layer1_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 8.705000 0.000000 8.845000 0.140000 ;
    END
  END start_layer1_i
  PIN start_layer2_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 10.665000 0.000000 10.805000 0.140000 ;
    END
  END start_layer2_i
  PIN weight_bias_mem_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 12.345000 0.000000 12.485000 0.140000 ;
    END
  END weight_bias_mem_req_o
  PIN weight_bias_mem_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 14.305000 0.000000 14.445000 0.140000 ;
    END
  END weight_bias_mem_ack_i
  PIN weight_bias_mem_addr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 72.825000 437.430000 72.965000 437.570000 ;
    END
  END weight_bias_mem_addr_o[9]
  PIN weight_bias_mem_addr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 73.665000 437.430000 73.805000 437.570000 ;
    END
  END weight_bias_mem_addr_o[8]
  PIN weight_bias_mem_addr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 74.505000 437.430000 74.645000 437.570000 ;
    END
  END weight_bias_mem_addr_o[7]
  PIN weight_bias_mem_addr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 75.345000 437.430000 75.485000 437.570000 ;
    END
  END weight_bias_mem_addr_o[6]
  PIN weight_bias_mem_addr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 76.185000 437.430000 76.325000 437.570000 ;
    END
  END weight_bias_mem_addr_o[5]
  PIN weight_bias_mem_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 77.025000 437.430000 77.165000 437.570000 ;
    END
  END weight_bias_mem_addr_o[4]
  PIN weight_bias_mem_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 77.865000 437.430000 78.005000 437.570000 ;
    END
  END weight_bias_mem_addr_o[3]
  PIN weight_bias_mem_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 78.705000 437.430000 78.845000 437.570000 ;
    END
  END weight_bias_mem_addr_o[2]
  PIN weight_bias_mem_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 79.545000 437.430000 79.685000 437.570000 ;
    END
  END weight_bias_mem_addr_o[1]
  PIN weight_bias_mem_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 80.385000 437.430000 80.525000 437.570000 ;
    END
  END weight_bias_mem_addr_o[0]
  PIN img_mem_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 16.265000 0.000000 16.405000 0.140000 ;
    END
  END img_mem_req_o
  PIN img_mem_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 17.945000 0.000000 18.085000 0.140000 ;
    END
  END img_mem_ack_i
  PIN img_mem_addr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 144.425000 0.140000 144.565000 ;
    END
  END img_mem_addr_o[4]
  PIN img_mem_addr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 144.995000 0.140000 145.135000 ;
    END
  END img_mem_addr_o[3]
  PIN img_mem_addr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 145.565000 0.140000 145.705000 ;
    END
  END img_mem_addr_o[2]
  PIN img_mem_addr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 146.135000 0.140000 146.275000 ;
    END
  END img_mem_addr_o[1]
  PIN img_mem_addr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 146.705000 0.140000 146.845000 ;
    END
  END img_mem_addr_o[0]
  PIN layer1_done_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 19.905000 0.000000 20.045000 0.140000 ;
    END
  END layer1_done_o
  PIN layer2_done_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 21.585000 0.000000 21.725000 0.140000 ;
    END
  END layer2_done_o
  PIN image_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 147.275000 0.140000 147.415000 ;
    END
  END image_i[255]
  PIN image_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 147.845000 0.140000 147.985000 ;
    END
  END image_i[254]
  PIN image_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 148.415000 0.140000 148.555000 ;
    END
  END image_i[253]
  PIN image_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 148.985000 0.140000 149.125000 ;
    END
  END image_i[252]
  PIN image_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 149.555000 0.140000 149.695000 ;
    END
  END image_i[251]
  PIN image_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 150.125000 0.140000 150.265000 ;
    END
  END image_i[250]
  PIN image_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 150.695000 0.140000 150.835000 ;
    END
  END image_i[249]
  PIN image_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 151.265000 0.140000 151.405000 ;
    END
  END image_i[248]
  PIN image_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 151.835000 0.140000 151.975000 ;
    END
  END image_i[247]
  PIN image_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 152.405000 0.140000 152.545000 ;
    END
  END image_i[246]
  PIN image_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 152.975000 0.140000 153.115000 ;
    END
  END image_i[245]
  PIN image_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 153.545000 0.140000 153.685000 ;
    END
  END image_i[244]
  PIN image_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 154.115000 0.140000 154.255000 ;
    END
  END image_i[243]
  PIN image_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 154.685000 0.140000 154.825000 ;
    END
  END image_i[242]
  PIN image_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 155.255000 0.140000 155.395000 ;
    END
  END image_i[241]
  PIN image_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 155.825000 0.140000 155.965000 ;
    END
  END image_i[240]
  PIN image_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 156.395000 0.140000 156.535000 ;
    END
  END image_i[239]
  PIN image_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 156.965000 0.140000 157.105000 ;
    END
  END image_i[238]
  PIN image_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 157.535000 0.140000 157.675000 ;
    END
  END image_i[237]
  PIN image_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 158.105000 0.140000 158.245000 ;
    END
  END image_i[236]
  PIN image_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 158.675000 0.140000 158.815000 ;
    END
  END image_i[235]
  PIN image_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 159.245000 0.140000 159.385000 ;
    END
  END image_i[234]
  PIN image_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 159.815000 0.140000 159.955000 ;
    END
  END image_i[233]
  PIN image_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 160.385000 0.140000 160.525000 ;
    END
  END image_i[232]
  PIN image_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 160.955000 0.140000 161.095000 ;
    END
  END image_i[231]
  PIN image_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 161.525000 0.140000 161.665000 ;
    END
  END image_i[230]
  PIN image_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 162.095000 0.140000 162.235000 ;
    END
  END image_i[229]
  PIN image_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 162.665000 0.140000 162.805000 ;
    END
  END image_i[228]
  PIN image_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 163.235000 0.140000 163.375000 ;
    END
  END image_i[227]
  PIN image_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 163.805000 0.140000 163.945000 ;
    END
  END image_i[226]
  PIN image_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 164.375000 0.140000 164.515000 ;
    END
  END image_i[225]
  PIN image_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 164.945000 0.140000 165.085000 ;
    END
  END image_i[224]
  PIN image_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 165.515000 0.140000 165.655000 ;
    END
  END image_i[223]
  PIN image_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 166.085000 0.140000 166.225000 ;
    END
  END image_i[222]
  PIN image_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 166.655000 0.140000 166.795000 ;
    END
  END image_i[221]
  PIN image_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 167.225000 0.140000 167.365000 ;
    END
  END image_i[220]
  PIN image_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 167.795000 0.140000 167.935000 ;
    END
  END image_i[219]
  PIN image_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 168.365000 0.140000 168.505000 ;
    END
  END image_i[218]
  PIN image_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 168.935000 0.140000 169.075000 ;
    END
  END image_i[217]
  PIN image_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 169.505000 0.140000 169.645000 ;
    END
  END image_i[216]
  PIN image_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 170.075000 0.140000 170.215000 ;
    END
  END image_i[215]
  PIN image_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 170.645000 0.140000 170.785000 ;
    END
  END image_i[214]
  PIN image_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 171.215000 0.140000 171.355000 ;
    END
  END image_i[213]
  PIN image_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 171.785000 0.140000 171.925000 ;
    END
  END image_i[212]
  PIN image_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 172.355000 0.140000 172.495000 ;
    END
  END image_i[211]
  PIN image_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 172.925000 0.140000 173.065000 ;
    END
  END image_i[210]
  PIN image_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 173.495000 0.140000 173.635000 ;
    END
  END image_i[209]
  PIN image_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 174.065000 0.140000 174.205000 ;
    END
  END image_i[208]
  PIN image_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 174.635000 0.140000 174.775000 ;
    END
  END image_i[207]
  PIN image_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 175.205000 0.140000 175.345000 ;
    END
  END image_i[206]
  PIN image_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 175.775000 0.140000 175.915000 ;
    END
  END image_i[205]
  PIN image_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 176.345000 0.140000 176.485000 ;
    END
  END image_i[204]
  PIN image_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 176.915000 0.140000 177.055000 ;
    END
  END image_i[203]
  PIN image_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 177.485000 0.140000 177.625000 ;
    END
  END image_i[202]
  PIN image_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 178.055000 0.140000 178.195000 ;
    END
  END image_i[201]
  PIN image_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 178.625000 0.140000 178.765000 ;
    END
  END image_i[200]
  PIN image_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 179.195000 0.140000 179.335000 ;
    END
  END image_i[199]
  PIN image_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 179.765000 0.140000 179.905000 ;
    END
  END image_i[198]
  PIN image_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 180.335000 0.140000 180.475000 ;
    END
  END image_i[197]
  PIN image_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 180.905000 0.140000 181.045000 ;
    END
  END image_i[196]
  PIN image_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 181.475000 0.140000 181.615000 ;
    END
  END image_i[195]
  PIN image_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 182.045000 0.140000 182.185000 ;
    END
  END image_i[194]
  PIN image_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 182.615000 0.140000 182.755000 ;
    END
  END image_i[193]
  PIN image_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 183.185000 0.140000 183.325000 ;
    END
  END image_i[192]
  PIN image_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 183.755000 0.140000 183.895000 ;
    END
  END image_i[191]
  PIN image_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 184.325000 0.140000 184.465000 ;
    END
  END image_i[190]
  PIN image_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 184.895000 0.140000 185.035000 ;
    END
  END image_i[189]
  PIN image_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 185.465000 0.140000 185.605000 ;
    END
  END image_i[188]
  PIN image_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 186.035000 0.140000 186.175000 ;
    END
  END image_i[187]
  PIN image_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 186.605000 0.140000 186.745000 ;
    END
  END image_i[186]
  PIN image_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 187.175000 0.140000 187.315000 ;
    END
  END image_i[185]
  PIN image_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 187.745000 0.140000 187.885000 ;
    END
  END image_i[184]
  PIN image_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 188.315000 0.140000 188.455000 ;
    END
  END image_i[183]
  PIN image_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 188.885000 0.140000 189.025000 ;
    END
  END image_i[182]
  PIN image_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 189.455000 0.140000 189.595000 ;
    END
  END image_i[181]
  PIN image_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 190.025000 0.140000 190.165000 ;
    END
  END image_i[180]
  PIN image_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 190.595000 0.140000 190.735000 ;
    END
  END image_i[179]
  PIN image_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 191.165000 0.140000 191.305000 ;
    END
  END image_i[178]
  PIN image_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 191.735000 0.140000 191.875000 ;
    END
  END image_i[177]
  PIN image_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 192.305000 0.140000 192.445000 ;
    END
  END image_i[176]
  PIN image_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 192.875000 0.140000 193.015000 ;
    END
  END image_i[175]
  PIN image_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 193.445000 0.140000 193.585000 ;
    END
  END image_i[174]
  PIN image_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 194.015000 0.140000 194.155000 ;
    END
  END image_i[173]
  PIN image_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 194.585000 0.140000 194.725000 ;
    END
  END image_i[172]
  PIN image_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 195.155000 0.140000 195.295000 ;
    END
  END image_i[171]
  PIN image_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 195.725000 0.140000 195.865000 ;
    END
  END image_i[170]
  PIN image_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 196.295000 0.140000 196.435000 ;
    END
  END image_i[169]
  PIN image_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 196.865000 0.140000 197.005000 ;
    END
  END image_i[168]
  PIN image_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 197.435000 0.140000 197.575000 ;
    END
  END image_i[167]
  PIN image_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 198.005000 0.140000 198.145000 ;
    END
  END image_i[166]
  PIN image_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 198.575000 0.140000 198.715000 ;
    END
  END image_i[165]
  PIN image_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 199.145000 0.140000 199.285000 ;
    END
  END image_i[164]
  PIN image_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 199.715000 0.140000 199.855000 ;
    END
  END image_i[163]
  PIN image_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 200.285000 0.140000 200.425000 ;
    END
  END image_i[162]
  PIN image_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 200.855000 0.140000 200.995000 ;
    END
  END image_i[161]
  PIN image_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 201.425000 0.140000 201.565000 ;
    END
  END image_i[160]
  PIN image_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 201.995000 0.140000 202.135000 ;
    END
  END image_i[159]
  PIN image_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 202.565000 0.140000 202.705000 ;
    END
  END image_i[158]
  PIN image_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 203.135000 0.140000 203.275000 ;
    END
  END image_i[157]
  PIN image_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 203.705000 0.140000 203.845000 ;
    END
  END image_i[156]
  PIN image_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 204.275000 0.140000 204.415000 ;
    END
  END image_i[155]
  PIN image_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 204.845000 0.140000 204.985000 ;
    END
  END image_i[154]
  PIN image_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 205.415000 0.140000 205.555000 ;
    END
  END image_i[153]
  PIN image_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 205.985000 0.140000 206.125000 ;
    END
  END image_i[152]
  PIN image_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 206.555000 0.140000 206.695000 ;
    END
  END image_i[151]
  PIN image_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 207.125000 0.140000 207.265000 ;
    END
  END image_i[150]
  PIN image_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 207.695000 0.140000 207.835000 ;
    END
  END image_i[149]
  PIN image_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 208.265000 0.140000 208.405000 ;
    END
  END image_i[148]
  PIN image_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 208.835000 0.140000 208.975000 ;
    END
  END image_i[147]
  PIN image_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 209.405000 0.140000 209.545000 ;
    END
  END image_i[146]
  PIN image_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 209.975000 0.140000 210.115000 ;
    END
  END image_i[145]
  PIN image_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 210.545000 0.140000 210.685000 ;
    END
  END image_i[144]
  PIN image_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 211.115000 0.140000 211.255000 ;
    END
  END image_i[143]
  PIN image_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 211.685000 0.140000 211.825000 ;
    END
  END image_i[142]
  PIN image_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 212.255000 0.140000 212.395000 ;
    END
  END image_i[141]
  PIN image_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 212.825000 0.140000 212.965000 ;
    END
  END image_i[140]
  PIN image_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 213.395000 0.140000 213.535000 ;
    END
  END image_i[139]
  PIN image_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 213.965000 0.140000 214.105000 ;
    END
  END image_i[138]
  PIN image_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 214.535000 0.140000 214.675000 ;
    END
  END image_i[137]
  PIN image_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 215.105000 0.140000 215.245000 ;
    END
  END image_i[136]
  PIN image_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 215.675000 0.140000 215.815000 ;
    END
  END image_i[135]
  PIN image_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 216.245000 0.140000 216.385000 ;
    END
  END image_i[134]
  PIN image_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 216.815000 0.140000 216.955000 ;
    END
  END image_i[133]
  PIN image_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 217.385000 0.140000 217.525000 ;
    END
  END image_i[132]
  PIN image_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 217.955000 0.140000 218.095000 ;
    END
  END image_i[131]
  PIN image_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 218.525000 0.140000 218.665000 ;
    END
  END image_i[130]
  PIN image_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 219.095000 0.140000 219.235000 ;
    END
  END image_i[129]
  PIN image_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 219.665000 0.140000 219.805000 ;
    END
  END image_i[128]
  PIN image_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 220.235000 0.140000 220.375000 ;
    END
  END image_i[127]
  PIN image_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 220.805000 0.140000 220.945000 ;
    END
  END image_i[126]
  PIN image_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 221.375000 0.140000 221.515000 ;
    END
  END image_i[125]
  PIN image_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 221.945000 0.140000 222.085000 ;
    END
  END image_i[124]
  PIN image_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 222.515000 0.140000 222.655000 ;
    END
  END image_i[123]
  PIN image_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 223.085000 0.140000 223.225000 ;
    END
  END image_i[122]
  PIN image_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 223.655000 0.140000 223.795000 ;
    END
  END image_i[121]
  PIN image_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 224.225000 0.140000 224.365000 ;
    END
  END image_i[120]
  PIN image_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 224.795000 0.140000 224.935000 ;
    END
  END image_i[119]
  PIN image_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 225.365000 0.140000 225.505000 ;
    END
  END image_i[118]
  PIN image_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 225.935000 0.140000 226.075000 ;
    END
  END image_i[117]
  PIN image_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 226.505000 0.140000 226.645000 ;
    END
  END image_i[116]
  PIN image_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 227.075000 0.140000 227.215000 ;
    END
  END image_i[115]
  PIN image_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 227.645000 0.140000 227.785000 ;
    END
  END image_i[114]
  PIN image_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 228.215000 0.140000 228.355000 ;
    END
  END image_i[113]
  PIN image_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 228.785000 0.140000 228.925000 ;
    END
  END image_i[112]
  PIN image_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 229.355000 0.140000 229.495000 ;
    END
  END image_i[111]
  PIN image_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 229.925000 0.140000 230.065000 ;
    END
  END image_i[110]
  PIN image_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 230.495000 0.140000 230.635000 ;
    END
  END image_i[109]
  PIN image_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 231.065000 0.140000 231.205000 ;
    END
  END image_i[108]
  PIN image_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 231.635000 0.140000 231.775000 ;
    END
  END image_i[107]
  PIN image_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 232.205000 0.140000 232.345000 ;
    END
  END image_i[106]
  PIN image_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 232.775000 0.140000 232.915000 ;
    END
  END image_i[105]
  PIN image_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 233.345000 0.140000 233.485000 ;
    END
  END image_i[104]
  PIN image_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 233.915000 0.140000 234.055000 ;
    END
  END image_i[103]
  PIN image_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 234.485000 0.140000 234.625000 ;
    END
  END image_i[102]
  PIN image_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 235.055000 0.140000 235.195000 ;
    END
  END image_i[101]
  PIN image_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 235.625000 0.140000 235.765000 ;
    END
  END image_i[100]
  PIN image_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 236.195000 0.140000 236.335000 ;
    END
  END image_i[99]
  PIN image_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 236.765000 0.140000 236.905000 ;
    END
  END image_i[98]
  PIN image_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 237.335000 0.140000 237.475000 ;
    END
  END image_i[97]
  PIN image_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 237.905000 0.140000 238.045000 ;
    END
  END image_i[96]
  PIN image_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 238.475000 0.140000 238.615000 ;
    END
  END image_i[95]
  PIN image_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 239.045000 0.140000 239.185000 ;
    END
  END image_i[94]
  PIN image_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 239.615000 0.140000 239.755000 ;
    END
  END image_i[93]
  PIN image_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 240.185000 0.140000 240.325000 ;
    END
  END image_i[92]
  PIN image_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 240.755000 0.140000 240.895000 ;
    END
  END image_i[91]
  PIN image_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 241.325000 0.140000 241.465000 ;
    END
  END image_i[90]
  PIN image_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 241.895000 0.140000 242.035000 ;
    END
  END image_i[89]
  PIN image_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 242.465000 0.140000 242.605000 ;
    END
  END image_i[88]
  PIN image_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 243.035000 0.140000 243.175000 ;
    END
  END image_i[87]
  PIN image_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 243.605000 0.140000 243.745000 ;
    END
  END image_i[86]
  PIN image_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 244.175000 0.140000 244.315000 ;
    END
  END image_i[85]
  PIN image_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 244.745000 0.140000 244.885000 ;
    END
  END image_i[84]
  PIN image_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 245.315000 0.140000 245.455000 ;
    END
  END image_i[83]
  PIN image_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 245.885000 0.140000 246.025000 ;
    END
  END image_i[82]
  PIN image_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 246.455000 0.140000 246.595000 ;
    END
  END image_i[81]
  PIN image_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 247.025000 0.140000 247.165000 ;
    END
  END image_i[80]
  PIN image_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 247.595000 0.140000 247.735000 ;
    END
  END image_i[79]
  PIN image_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 248.165000 0.140000 248.305000 ;
    END
  END image_i[78]
  PIN image_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 248.735000 0.140000 248.875000 ;
    END
  END image_i[77]
  PIN image_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 249.305000 0.140000 249.445000 ;
    END
  END image_i[76]
  PIN image_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 249.875000 0.140000 250.015000 ;
    END
  END image_i[75]
  PIN image_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 250.445000 0.140000 250.585000 ;
    END
  END image_i[74]
  PIN image_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 251.015000 0.140000 251.155000 ;
    END
  END image_i[73]
  PIN image_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 251.585000 0.140000 251.725000 ;
    END
  END image_i[72]
  PIN image_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 252.155000 0.140000 252.295000 ;
    END
  END image_i[71]
  PIN image_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 252.725000 0.140000 252.865000 ;
    END
  END image_i[70]
  PIN image_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 253.295000 0.140000 253.435000 ;
    END
  END image_i[69]
  PIN image_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 253.865000 0.140000 254.005000 ;
    END
  END image_i[68]
  PIN image_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 254.435000 0.140000 254.575000 ;
    END
  END image_i[67]
  PIN image_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 255.005000 0.140000 255.145000 ;
    END
  END image_i[66]
  PIN image_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 255.575000 0.140000 255.715000 ;
    END
  END image_i[65]
  PIN image_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 256.145000 0.140000 256.285000 ;
    END
  END image_i[64]
  PIN image_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 256.715000 0.140000 256.855000 ;
    END
  END image_i[63]
  PIN image_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 257.285000 0.140000 257.425000 ;
    END
  END image_i[62]
  PIN image_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 257.855000 0.140000 257.995000 ;
    END
  END image_i[61]
  PIN image_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 258.425000 0.140000 258.565000 ;
    END
  END image_i[60]
  PIN image_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 258.995000 0.140000 259.135000 ;
    END
  END image_i[59]
  PIN image_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 259.565000 0.140000 259.705000 ;
    END
  END image_i[58]
  PIN image_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 260.135000 0.140000 260.275000 ;
    END
  END image_i[57]
  PIN image_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 260.705000 0.140000 260.845000 ;
    END
  END image_i[56]
  PIN image_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 261.275000 0.140000 261.415000 ;
    END
  END image_i[55]
  PIN image_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 261.845000 0.140000 261.985000 ;
    END
  END image_i[54]
  PIN image_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 262.415000 0.140000 262.555000 ;
    END
  END image_i[53]
  PIN image_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 262.985000 0.140000 263.125000 ;
    END
  END image_i[52]
  PIN image_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 263.555000 0.140000 263.695000 ;
    END
  END image_i[51]
  PIN image_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 264.125000 0.140000 264.265000 ;
    END
  END image_i[50]
  PIN image_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 264.695000 0.140000 264.835000 ;
    END
  END image_i[49]
  PIN image_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 265.265000 0.140000 265.405000 ;
    END
  END image_i[48]
  PIN image_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 265.835000 0.140000 265.975000 ;
    END
  END image_i[47]
  PIN image_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 266.405000 0.140000 266.545000 ;
    END
  END image_i[46]
  PIN image_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 266.975000 0.140000 267.115000 ;
    END
  END image_i[45]
  PIN image_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 267.545000 0.140000 267.685000 ;
    END
  END image_i[44]
  PIN image_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 268.115000 0.140000 268.255000 ;
    END
  END image_i[43]
  PIN image_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 268.685000 0.140000 268.825000 ;
    END
  END image_i[42]
  PIN image_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 269.255000 0.140000 269.395000 ;
    END
  END image_i[41]
  PIN image_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 269.825000 0.140000 269.965000 ;
    END
  END image_i[40]
  PIN image_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 270.395000 0.140000 270.535000 ;
    END
  END image_i[39]
  PIN image_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 270.965000 0.140000 271.105000 ;
    END
  END image_i[38]
  PIN image_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 271.535000 0.140000 271.675000 ;
    END
  END image_i[37]
  PIN image_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 272.105000 0.140000 272.245000 ;
    END
  END image_i[36]
  PIN image_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 272.675000 0.140000 272.815000 ;
    END
  END image_i[35]
  PIN image_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 273.245000 0.140000 273.385000 ;
    END
  END image_i[34]
  PIN image_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 273.815000 0.140000 273.955000 ;
    END
  END image_i[33]
  PIN image_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 274.385000 0.140000 274.525000 ;
    END
  END image_i[32]
  PIN image_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 274.955000 0.140000 275.095000 ;
    END
  END image_i[31]
  PIN image_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 275.525000 0.140000 275.665000 ;
    END
  END image_i[30]
  PIN image_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 276.095000 0.140000 276.235000 ;
    END
  END image_i[29]
  PIN image_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 276.665000 0.140000 276.805000 ;
    END
  END image_i[28]
  PIN image_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 277.235000 0.140000 277.375000 ;
    END
  END image_i[27]
  PIN image_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 277.805000 0.140000 277.945000 ;
    END
  END image_i[26]
  PIN image_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 278.375000 0.140000 278.515000 ;
    END
  END image_i[25]
  PIN image_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 278.945000 0.140000 279.085000 ;
    END
  END image_i[24]
  PIN image_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 279.515000 0.140000 279.655000 ;
    END
  END image_i[23]
  PIN image_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 280.085000 0.140000 280.225000 ;
    END
  END image_i[22]
  PIN image_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 280.655000 0.140000 280.795000 ;
    END
  END image_i[21]
  PIN image_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 281.225000 0.140000 281.365000 ;
    END
  END image_i[20]
  PIN image_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 281.795000 0.140000 281.935000 ;
    END
  END image_i[19]
  PIN image_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 282.365000 0.140000 282.505000 ;
    END
  END image_i[18]
  PIN image_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 282.935000 0.140000 283.075000 ;
    END
  END image_i[17]
  PIN image_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 283.505000 0.140000 283.645000 ;
    END
  END image_i[16]
  PIN image_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 284.075000 0.140000 284.215000 ;
    END
  END image_i[15]
  PIN image_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 284.645000 0.140000 284.785000 ;
    END
  END image_i[14]
  PIN image_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 285.215000 0.140000 285.355000 ;
    END
  END image_i[13]
  PIN image_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 285.785000 0.140000 285.925000 ;
    END
  END image_i[12]
  PIN image_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 286.355000 0.140000 286.495000 ;
    END
  END image_i[11]
  PIN image_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 286.925000 0.140000 287.065000 ;
    END
  END image_i[10]
  PIN image_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 287.495000 0.140000 287.635000 ;
    END
  END image_i[9]
  PIN image_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 288.065000 0.140000 288.205000 ;
    END
  END image_i[8]
  PIN image_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 288.635000 0.140000 288.775000 ;
    END
  END image_i[7]
  PIN image_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 289.205000 0.140000 289.345000 ;
    END
  END image_i[6]
  PIN image_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 289.775000 0.140000 289.915000 ;
    END
  END image_i[5]
  PIN image_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 290.345000 0.140000 290.485000 ;
    END
  END image_i[4]
  PIN image_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 290.915000 0.140000 291.055000 ;
    END
  END image_i[3]
  PIN image_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 291.485000 0.140000 291.625000 ;
    END
  END image_i[2]
  PIN image_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 292.055000 0.140000 292.195000 ;
    END
  END image_i[1]
  PIN image_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 0.000000 292.625000 0.140000 292.765000 ;
    END
  END image_i[0]
  PIN weight_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 81.225000 437.430000 81.365000 437.570000 ;
    END
  END weight_i[255]
  PIN weight_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 82.065000 437.430000 82.205000 437.570000 ;
    END
  END weight_i[254]
  PIN weight_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 82.905000 437.430000 83.045000 437.570000 ;
    END
  END weight_i[253]
  PIN weight_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 83.745000 437.430000 83.885000 437.570000 ;
    END
  END weight_i[252]
  PIN weight_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 84.585000 437.430000 84.725000 437.570000 ;
    END
  END weight_i[251]
  PIN weight_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 85.425000 437.430000 85.565000 437.570000 ;
    END
  END weight_i[250]
  PIN weight_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 86.265000 437.430000 86.405000 437.570000 ;
    END
  END weight_i[249]
  PIN weight_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 87.105000 437.430000 87.245000 437.570000 ;
    END
  END weight_i[248]
  PIN weight_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 87.945000 437.430000 88.085000 437.570000 ;
    END
  END weight_i[247]
  PIN weight_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 88.785000 437.430000 88.925000 437.570000 ;
    END
  END weight_i[246]
  PIN weight_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 89.625000 437.430000 89.765000 437.570000 ;
    END
  END weight_i[245]
  PIN weight_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 90.465000 437.430000 90.605000 437.570000 ;
    END
  END weight_i[244]
  PIN weight_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 91.305000 437.430000 91.445000 437.570000 ;
    END
  END weight_i[243]
  PIN weight_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 92.145000 437.430000 92.285000 437.570000 ;
    END
  END weight_i[242]
  PIN weight_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 92.985000 437.430000 93.125000 437.570000 ;
    END
  END weight_i[241]
  PIN weight_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 93.825000 437.430000 93.965000 437.570000 ;
    END
  END weight_i[240]
  PIN weight_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 94.665000 437.430000 94.805000 437.570000 ;
    END
  END weight_i[239]
  PIN weight_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 95.505000 437.430000 95.645000 437.570000 ;
    END
  END weight_i[238]
  PIN weight_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 96.345000 437.430000 96.485000 437.570000 ;
    END
  END weight_i[237]
  PIN weight_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 97.185000 437.430000 97.325000 437.570000 ;
    END
  END weight_i[236]
  PIN weight_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 98.025000 437.430000 98.165000 437.570000 ;
    END
  END weight_i[235]
  PIN weight_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 98.865000 437.430000 99.005000 437.570000 ;
    END
  END weight_i[234]
  PIN weight_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 99.705000 437.430000 99.845000 437.570000 ;
    END
  END weight_i[233]
  PIN weight_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 100.545000 437.430000 100.685000 437.570000 ;
    END
  END weight_i[232]
  PIN weight_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 101.385000 437.430000 101.525000 437.570000 ;
    END
  END weight_i[231]
  PIN weight_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 102.225000 437.430000 102.365000 437.570000 ;
    END
  END weight_i[230]
  PIN weight_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 103.065000 437.430000 103.205000 437.570000 ;
    END
  END weight_i[229]
  PIN weight_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 103.905000 437.430000 104.045000 437.570000 ;
    END
  END weight_i[228]
  PIN weight_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 104.745000 437.430000 104.885000 437.570000 ;
    END
  END weight_i[227]
  PIN weight_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 105.585000 437.430000 105.725000 437.570000 ;
    END
  END weight_i[226]
  PIN weight_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 106.425000 437.430000 106.565000 437.570000 ;
    END
  END weight_i[225]
  PIN weight_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 107.265000 437.430000 107.405000 437.570000 ;
    END
  END weight_i[224]
  PIN weight_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 108.105000 437.430000 108.245000 437.570000 ;
    END
  END weight_i[223]
  PIN weight_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 108.945000 437.430000 109.085000 437.570000 ;
    END
  END weight_i[222]
  PIN weight_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 109.785000 437.430000 109.925000 437.570000 ;
    END
  END weight_i[221]
  PIN weight_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 110.625000 437.430000 110.765000 437.570000 ;
    END
  END weight_i[220]
  PIN weight_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 111.465000 437.430000 111.605000 437.570000 ;
    END
  END weight_i[219]
  PIN weight_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 112.305000 437.430000 112.445000 437.570000 ;
    END
  END weight_i[218]
  PIN weight_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 113.145000 437.430000 113.285000 437.570000 ;
    END
  END weight_i[217]
  PIN weight_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 113.985000 437.430000 114.125000 437.570000 ;
    END
  END weight_i[216]
  PIN weight_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 114.825000 437.430000 114.965000 437.570000 ;
    END
  END weight_i[215]
  PIN weight_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 115.665000 437.430000 115.805000 437.570000 ;
    END
  END weight_i[214]
  PIN weight_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 116.505000 437.430000 116.645000 437.570000 ;
    END
  END weight_i[213]
  PIN weight_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 117.345000 437.430000 117.485000 437.570000 ;
    END
  END weight_i[212]
  PIN weight_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 118.185000 437.430000 118.325000 437.570000 ;
    END
  END weight_i[211]
  PIN weight_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 119.025000 437.430000 119.165000 437.570000 ;
    END
  END weight_i[210]
  PIN weight_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 119.865000 437.430000 120.005000 437.570000 ;
    END
  END weight_i[209]
  PIN weight_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 120.705000 437.430000 120.845000 437.570000 ;
    END
  END weight_i[208]
  PIN weight_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 121.545000 437.430000 121.685000 437.570000 ;
    END
  END weight_i[207]
  PIN weight_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 122.385000 437.430000 122.525000 437.570000 ;
    END
  END weight_i[206]
  PIN weight_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 123.225000 437.430000 123.365000 437.570000 ;
    END
  END weight_i[205]
  PIN weight_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 124.065000 437.430000 124.205000 437.570000 ;
    END
  END weight_i[204]
  PIN weight_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 124.905000 437.430000 125.045000 437.570000 ;
    END
  END weight_i[203]
  PIN weight_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 125.745000 437.430000 125.885000 437.570000 ;
    END
  END weight_i[202]
  PIN weight_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 126.585000 437.430000 126.725000 437.570000 ;
    END
  END weight_i[201]
  PIN weight_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 127.425000 437.430000 127.565000 437.570000 ;
    END
  END weight_i[200]
  PIN weight_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 128.265000 437.430000 128.405000 437.570000 ;
    END
  END weight_i[199]
  PIN weight_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 129.105000 437.430000 129.245000 437.570000 ;
    END
  END weight_i[198]
  PIN weight_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 129.945000 437.430000 130.085000 437.570000 ;
    END
  END weight_i[197]
  PIN weight_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 130.785000 437.430000 130.925000 437.570000 ;
    END
  END weight_i[196]
  PIN weight_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 131.625000 437.430000 131.765000 437.570000 ;
    END
  END weight_i[195]
  PIN weight_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 132.465000 437.430000 132.605000 437.570000 ;
    END
  END weight_i[194]
  PIN weight_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 133.305000 437.430000 133.445000 437.570000 ;
    END
  END weight_i[193]
  PIN weight_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 134.145000 437.430000 134.285000 437.570000 ;
    END
  END weight_i[192]
  PIN weight_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 134.985000 437.430000 135.125000 437.570000 ;
    END
  END weight_i[191]
  PIN weight_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 135.825000 437.430000 135.965000 437.570000 ;
    END
  END weight_i[190]
  PIN weight_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 136.665000 437.430000 136.805000 437.570000 ;
    END
  END weight_i[189]
  PIN weight_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 137.505000 437.430000 137.645000 437.570000 ;
    END
  END weight_i[188]
  PIN weight_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 138.345000 437.430000 138.485000 437.570000 ;
    END
  END weight_i[187]
  PIN weight_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 139.185000 437.430000 139.325000 437.570000 ;
    END
  END weight_i[186]
  PIN weight_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 140.025000 437.430000 140.165000 437.570000 ;
    END
  END weight_i[185]
  PIN weight_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 140.865000 437.430000 141.005000 437.570000 ;
    END
  END weight_i[184]
  PIN weight_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 141.705000 437.430000 141.845000 437.570000 ;
    END
  END weight_i[183]
  PIN weight_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 142.545000 437.430000 142.685000 437.570000 ;
    END
  END weight_i[182]
  PIN weight_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 143.385000 437.430000 143.525000 437.570000 ;
    END
  END weight_i[181]
  PIN weight_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 144.225000 437.430000 144.365000 437.570000 ;
    END
  END weight_i[180]
  PIN weight_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 145.065000 437.430000 145.205000 437.570000 ;
    END
  END weight_i[179]
  PIN weight_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 145.905000 437.430000 146.045000 437.570000 ;
    END
  END weight_i[178]
  PIN weight_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 146.745000 437.430000 146.885000 437.570000 ;
    END
  END weight_i[177]
  PIN weight_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 147.585000 437.430000 147.725000 437.570000 ;
    END
  END weight_i[176]
  PIN weight_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 148.425000 437.430000 148.565000 437.570000 ;
    END
  END weight_i[175]
  PIN weight_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 149.265000 437.430000 149.405000 437.570000 ;
    END
  END weight_i[174]
  PIN weight_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 150.105000 437.430000 150.245000 437.570000 ;
    END
  END weight_i[173]
  PIN weight_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 150.945000 437.430000 151.085000 437.570000 ;
    END
  END weight_i[172]
  PIN weight_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 151.785000 437.430000 151.925000 437.570000 ;
    END
  END weight_i[171]
  PIN weight_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 152.625000 437.430000 152.765000 437.570000 ;
    END
  END weight_i[170]
  PIN weight_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 153.465000 437.430000 153.605000 437.570000 ;
    END
  END weight_i[169]
  PIN weight_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 154.305000 437.430000 154.445000 437.570000 ;
    END
  END weight_i[168]
  PIN weight_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 155.145000 437.430000 155.285000 437.570000 ;
    END
  END weight_i[167]
  PIN weight_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 155.985000 437.430000 156.125000 437.570000 ;
    END
  END weight_i[166]
  PIN weight_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 156.825000 437.430000 156.965000 437.570000 ;
    END
  END weight_i[165]
  PIN weight_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 157.665000 437.430000 157.805000 437.570000 ;
    END
  END weight_i[164]
  PIN weight_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 158.505000 437.430000 158.645000 437.570000 ;
    END
  END weight_i[163]
  PIN weight_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 159.345000 437.430000 159.485000 437.570000 ;
    END
  END weight_i[162]
  PIN weight_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 160.185000 437.430000 160.325000 437.570000 ;
    END
  END weight_i[161]
  PIN weight_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 161.025000 437.430000 161.165000 437.570000 ;
    END
  END weight_i[160]
  PIN weight_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 161.865000 437.430000 162.005000 437.570000 ;
    END
  END weight_i[159]
  PIN weight_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 162.705000 437.430000 162.845000 437.570000 ;
    END
  END weight_i[158]
  PIN weight_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 163.545000 437.430000 163.685000 437.570000 ;
    END
  END weight_i[157]
  PIN weight_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 164.385000 437.430000 164.525000 437.570000 ;
    END
  END weight_i[156]
  PIN weight_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 165.225000 437.430000 165.365000 437.570000 ;
    END
  END weight_i[155]
  PIN weight_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 166.065000 437.430000 166.205000 437.570000 ;
    END
  END weight_i[154]
  PIN weight_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 166.905000 437.430000 167.045000 437.570000 ;
    END
  END weight_i[153]
  PIN weight_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 167.745000 437.430000 167.885000 437.570000 ;
    END
  END weight_i[152]
  PIN weight_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 168.585000 437.430000 168.725000 437.570000 ;
    END
  END weight_i[151]
  PIN weight_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 169.425000 437.430000 169.565000 437.570000 ;
    END
  END weight_i[150]
  PIN weight_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 170.265000 437.430000 170.405000 437.570000 ;
    END
  END weight_i[149]
  PIN weight_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 171.105000 437.430000 171.245000 437.570000 ;
    END
  END weight_i[148]
  PIN weight_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 171.945000 437.430000 172.085000 437.570000 ;
    END
  END weight_i[147]
  PIN weight_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 172.785000 437.430000 172.925000 437.570000 ;
    END
  END weight_i[146]
  PIN weight_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 173.625000 437.430000 173.765000 437.570000 ;
    END
  END weight_i[145]
  PIN weight_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 174.465000 437.430000 174.605000 437.570000 ;
    END
  END weight_i[144]
  PIN weight_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 175.305000 437.430000 175.445000 437.570000 ;
    END
  END weight_i[143]
  PIN weight_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 176.145000 437.430000 176.285000 437.570000 ;
    END
  END weight_i[142]
  PIN weight_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 176.985000 437.430000 177.125000 437.570000 ;
    END
  END weight_i[141]
  PIN weight_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 177.825000 437.430000 177.965000 437.570000 ;
    END
  END weight_i[140]
  PIN weight_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 178.665000 437.430000 178.805000 437.570000 ;
    END
  END weight_i[139]
  PIN weight_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 179.505000 437.430000 179.645000 437.570000 ;
    END
  END weight_i[138]
  PIN weight_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 180.345000 437.430000 180.485000 437.570000 ;
    END
  END weight_i[137]
  PIN weight_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 181.185000 437.430000 181.325000 437.570000 ;
    END
  END weight_i[136]
  PIN weight_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 182.025000 437.430000 182.165000 437.570000 ;
    END
  END weight_i[135]
  PIN weight_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 182.865000 437.430000 183.005000 437.570000 ;
    END
  END weight_i[134]
  PIN weight_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 183.705000 437.430000 183.845000 437.570000 ;
    END
  END weight_i[133]
  PIN weight_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 184.545000 437.430000 184.685000 437.570000 ;
    END
  END weight_i[132]
  PIN weight_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 185.385000 437.430000 185.525000 437.570000 ;
    END
  END weight_i[131]
  PIN weight_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 186.225000 437.430000 186.365000 437.570000 ;
    END
  END weight_i[130]
  PIN weight_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 187.065000 437.430000 187.205000 437.570000 ;
    END
  END weight_i[129]
  PIN weight_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 187.905000 437.430000 188.045000 437.570000 ;
    END
  END weight_i[128]
  PIN weight_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 188.745000 437.430000 188.885000 437.570000 ;
    END
  END weight_i[127]
  PIN weight_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 189.585000 437.430000 189.725000 437.570000 ;
    END
  END weight_i[126]
  PIN weight_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 190.425000 437.430000 190.565000 437.570000 ;
    END
  END weight_i[125]
  PIN weight_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 191.265000 437.430000 191.405000 437.570000 ;
    END
  END weight_i[124]
  PIN weight_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 192.105000 437.430000 192.245000 437.570000 ;
    END
  END weight_i[123]
  PIN weight_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 192.945000 437.430000 193.085000 437.570000 ;
    END
  END weight_i[122]
  PIN weight_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 193.785000 437.430000 193.925000 437.570000 ;
    END
  END weight_i[121]
  PIN weight_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 194.625000 437.430000 194.765000 437.570000 ;
    END
  END weight_i[120]
  PIN weight_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 195.465000 437.430000 195.605000 437.570000 ;
    END
  END weight_i[119]
  PIN weight_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 196.305000 437.430000 196.445000 437.570000 ;
    END
  END weight_i[118]
  PIN weight_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 197.145000 437.430000 197.285000 437.570000 ;
    END
  END weight_i[117]
  PIN weight_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 197.985000 437.430000 198.125000 437.570000 ;
    END
  END weight_i[116]
  PIN weight_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 198.825000 437.430000 198.965000 437.570000 ;
    END
  END weight_i[115]
  PIN weight_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 199.665000 437.430000 199.805000 437.570000 ;
    END
  END weight_i[114]
  PIN weight_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 200.505000 437.430000 200.645000 437.570000 ;
    END
  END weight_i[113]
  PIN weight_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 201.345000 437.430000 201.485000 437.570000 ;
    END
  END weight_i[112]
  PIN weight_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 202.185000 437.430000 202.325000 437.570000 ;
    END
  END weight_i[111]
  PIN weight_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 203.025000 437.430000 203.165000 437.570000 ;
    END
  END weight_i[110]
  PIN weight_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 203.865000 437.430000 204.005000 437.570000 ;
    END
  END weight_i[109]
  PIN weight_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 204.705000 437.430000 204.845000 437.570000 ;
    END
  END weight_i[108]
  PIN weight_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 205.545000 437.430000 205.685000 437.570000 ;
    END
  END weight_i[107]
  PIN weight_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 206.385000 437.430000 206.525000 437.570000 ;
    END
  END weight_i[106]
  PIN weight_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 207.225000 437.430000 207.365000 437.570000 ;
    END
  END weight_i[105]
  PIN weight_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 208.065000 437.430000 208.205000 437.570000 ;
    END
  END weight_i[104]
  PIN weight_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 208.905000 437.430000 209.045000 437.570000 ;
    END
  END weight_i[103]
  PIN weight_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 209.745000 437.430000 209.885000 437.570000 ;
    END
  END weight_i[102]
  PIN weight_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 210.585000 437.430000 210.725000 437.570000 ;
    END
  END weight_i[101]
  PIN weight_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 211.425000 437.430000 211.565000 437.570000 ;
    END
  END weight_i[100]
  PIN weight_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 212.265000 437.430000 212.405000 437.570000 ;
    END
  END weight_i[99]
  PIN weight_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 213.105000 437.430000 213.245000 437.570000 ;
    END
  END weight_i[98]
  PIN weight_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 213.945000 437.430000 214.085000 437.570000 ;
    END
  END weight_i[97]
  PIN weight_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 214.785000 437.430000 214.925000 437.570000 ;
    END
  END weight_i[96]
  PIN weight_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 215.625000 437.430000 215.765000 437.570000 ;
    END
  END weight_i[95]
  PIN weight_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 216.465000 437.430000 216.605000 437.570000 ;
    END
  END weight_i[94]
  PIN weight_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 217.305000 437.430000 217.445000 437.570000 ;
    END
  END weight_i[93]
  PIN weight_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 218.145000 437.430000 218.285000 437.570000 ;
    END
  END weight_i[92]
  PIN weight_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 218.985000 437.430000 219.125000 437.570000 ;
    END
  END weight_i[91]
  PIN weight_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 219.825000 437.430000 219.965000 437.570000 ;
    END
  END weight_i[90]
  PIN weight_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 220.665000 437.430000 220.805000 437.570000 ;
    END
  END weight_i[89]
  PIN weight_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 221.505000 437.430000 221.645000 437.570000 ;
    END
  END weight_i[88]
  PIN weight_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 222.345000 437.430000 222.485000 437.570000 ;
    END
  END weight_i[87]
  PIN weight_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 223.185000 437.430000 223.325000 437.570000 ;
    END
  END weight_i[86]
  PIN weight_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 224.025000 437.430000 224.165000 437.570000 ;
    END
  END weight_i[85]
  PIN weight_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 224.865000 437.430000 225.005000 437.570000 ;
    END
  END weight_i[84]
  PIN weight_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 225.705000 437.430000 225.845000 437.570000 ;
    END
  END weight_i[83]
  PIN weight_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 226.545000 437.430000 226.685000 437.570000 ;
    END
  END weight_i[82]
  PIN weight_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 227.385000 437.430000 227.525000 437.570000 ;
    END
  END weight_i[81]
  PIN weight_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 228.225000 437.430000 228.365000 437.570000 ;
    END
  END weight_i[80]
  PIN weight_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 229.065000 437.430000 229.205000 437.570000 ;
    END
  END weight_i[79]
  PIN weight_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 229.905000 437.430000 230.045000 437.570000 ;
    END
  END weight_i[78]
  PIN weight_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 230.745000 437.430000 230.885000 437.570000 ;
    END
  END weight_i[77]
  PIN weight_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 231.585000 437.430000 231.725000 437.570000 ;
    END
  END weight_i[76]
  PIN weight_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 232.425000 437.430000 232.565000 437.570000 ;
    END
  END weight_i[75]
  PIN weight_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 233.265000 437.430000 233.405000 437.570000 ;
    END
  END weight_i[74]
  PIN weight_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 234.105000 437.430000 234.245000 437.570000 ;
    END
  END weight_i[73]
  PIN weight_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 234.945000 437.430000 235.085000 437.570000 ;
    END
  END weight_i[72]
  PIN weight_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 235.785000 437.430000 235.925000 437.570000 ;
    END
  END weight_i[71]
  PIN weight_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 236.625000 437.430000 236.765000 437.570000 ;
    END
  END weight_i[70]
  PIN weight_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 237.465000 437.430000 237.605000 437.570000 ;
    END
  END weight_i[69]
  PIN weight_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 238.305000 437.430000 238.445000 437.570000 ;
    END
  END weight_i[68]
  PIN weight_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 239.145000 437.430000 239.285000 437.570000 ;
    END
  END weight_i[67]
  PIN weight_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 239.985000 437.430000 240.125000 437.570000 ;
    END
  END weight_i[66]
  PIN weight_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 240.825000 437.430000 240.965000 437.570000 ;
    END
  END weight_i[65]
  PIN weight_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 241.665000 437.430000 241.805000 437.570000 ;
    END
  END weight_i[64]
  PIN weight_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 242.505000 437.430000 242.645000 437.570000 ;
    END
  END weight_i[63]
  PIN weight_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 243.345000 437.430000 243.485000 437.570000 ;
    END
  END weight_i[62]
  PIN weight_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 244.185000 437.430000 244.325000 437.570000 ;
    END
  END weight_i[61]
  PIN weight_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 245.025000 437.430000 245.165000 437.570000 ;
    END
  END weight_i[60]
  PIN weight_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 245.865000 437.430000 246.005000 437.570000 ;
    END
  END weight_i[59]
  PIN weight_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 246.705000 437.430000 246.845000 437.570000 ;
    END
  END weight_i[58]
  PIN weight_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 247.545000 437.430000 247.685000 437.570000 ;
    END
  END weight_i[57]
  PIN weight_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 248.385000 437.430000 248.525000 437.570000 ;
    END
  END weight_i[56]
  PIN weight_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 249.225000 437.430000 249.365000 437.570000 ;
    END
  END weight_i[55]
  PIN weight_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 250.065000 437.430000 250.205000 437.570000 ;
    END
  END weight_i[54]
  PIN weight_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 250.905000 437.430000 251.045000 437.570000 ;
    END
  END weight_i[53]
  PIN weight_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 251.745000 437.430000 251.885000 437.570000 ;
    END
  END weight_i[52]
  PIN weight_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 252.585000 437.430000 252.725000 437.570000 ;
    END
  END weight_i[51]
  PIN weight_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 253.425000 437.430000 253.565000 437.570000 ;
    END
  END weight_i[50]
  PIN weight_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 254.265000 437.430000 254.405000 437.570000 ;
    END
  END weight_i[49]
  PIN weight_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 255.105000 437.430000 255.245000 437.570000 ;
    END
  END weight_i[48]
  PIN weight_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 255.945000 437.430000 256.085000 437.570000 ;
    END
  END weight_i[47]
  PIN weight_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 256.785000 437.430000 256.925000 437.570000 ;
    END
  END weight_i[46]
  PIN weight_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 257.625000 437.430000 257.765000 437.570000 ;
    END
  END weight_i[45]
  PIN weight_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 258.465000 437.430000 258.605000 437.570000 ;
    END
  END weight_i[44]
  PIN weight_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 259.305000 437.430000 259.445000 437.570000 ;
    END
  END weight_i[43]
  PIN weight_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 260.145000 437.430000 260.285000 437.570000 ;
    END
  END weight_i[42]
  PIN weight_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 260.985000 437.430000 261.125000 437.570000 ;
    END
  END weight_i[41]
  PIN weight_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 261.825000 437.430000 261.965000 437.570000 ;
    END
  END weight_i[40]
  PIN weight_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 262.665000 437.430000 262.805000 437.570000 ;
    END
  END weight_i[39]
  PIN weight_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 263.505000 437.430000 263.645000 437.570000 ;
    END
  END weight_i[38]
  PIN weight_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 264.345000 437.430000 264.485000 437.570000 ;
    END
  END weight_i[37]
  PIN weight_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 265.185000 437.430000 265.325000 437.570000 ;
    END
  END weight_i[36]
  PIN weight_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 266.025000 437.430000 266.165000 437.570000 ;
    END
  END weight_i[35]
  PIN weight_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 266.865000 437.430000 267.005000 437.570000 ;
    END
  END weight_i[34]
  PIN weight_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 267.705000 437.430000 267.845000 437.570000 ;
    END
  END weight_i[33]
  PIN weight_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 268.545000 437.430000 268.685000 437.570000 ;
    END
  END weight_i[32]
  PIN weight_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 269.385000 437.430000 269.525000 437.570000 ;
    END
  END weight_i[31]
  PIN weight_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 270.225000 437.430000 270.365000 437.570000 ;
    END
  END weight_i[30]
  PIN weight_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 271.065000 437.430000 271.205000 437.570000 ;
    END
  END weight_i[29]
  PIN weight_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 271.905000 437.430000 272.045000 437.570000 ;
    END
  END weight_i[28]
  PIN weight_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 272.745000 437.430000 272.885000 437.570000 ;
    END
  END weight_i[27]
  PIN weight_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 273.585000 437.430000 273.725000 437.570000 ;
    END
  END weight_i[26]
  PIN weight_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 274.425000 437.430000 274.565000 437.570000 ;
    END
  END weight_i[25]
  PIN weight_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 275.265000 437.430000 275.405000 437.570000 ;
    END
  END weight_i[24]
  PIN weight_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 276.105000 437.430000 276.245000 437.570000 ;
    END
  END weight_i[23]
  PIN weight_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 276.945000 437.430000 277.085000 437.570000 ;
    END
  END weight_i[22]
  PIN weight_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 277.785000 437.430000 277.925000 437.570000 ;
    END
  END weight_i[21]
  PIN weight_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 278.625000 437.430000 278.765000 437.570000 ;
    END
  END weight_i[20]
  PIN weight_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 279.465000 437.430000 279.605000 437.570000 ;
    END
  END weight_i[19]
  PIN weight_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 280.305000 437.430000 280.445000 437.570000 ;
    END
  END weight_i[18]
  PIN weight_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 281.145000 437.430000 281.285000 437.570000 ;
    END
  END weight_i[17]
  PIN weight_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 281.985000 437.430000 282.125000 437.570000 ;
    END
  END weight_i[16]
  PIN weight_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 282.825000 437.430000 282.965000 437.570000 ;
    END
  END weight_i[15]
  PIN weight_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 283.665000 437.430000 283.805000 437.570000 ;
    END
  END weight_i[14]
  PIN weight_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 284.505000 437.430000 284.645000 437.570000 ;
    END
  END weight_i[13]
  PIN weight_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 285.345000 437.430000 285.485000 437.570000 ;
    END
  END weight_i[12]
  PIN weight_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 286.185000 437.430000 286.325000 437.570000 ;
    END
  END weight_i[11]
  PIN weight_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 287.025000 437.430000 287.165000 437.570000 ;
    END
  END weight_i[10]
  PIN weight_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 287.865000 437.430000 288.005000 437.570000 ;
    END
  END weight_i[9]
  PIN weight_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 288.705000 437.430000 288.845000 437.570000 ;
    END
  END weight_i[8]
  PIN weight_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 289.545000 437.430000 289.685000 437.570000 ;
    END
  END weight_i[7]
  PIN weight_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 290.385000 437.430000 290.525000 437.570000 ;
    END
  END weight_i[6]
  PIN weight_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 291.225000 437.430000 291.365000 437.570000 ;
    END
  END weight_i[5]
  PIN weight_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 292.065000 437.430000 292.205000 437.570000 ;
    END
  END weight_i[4]
  PIN weight_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 292.905000 437.430000 293.045000 437.570000 ;
    END
  END weight_i[3]
  PIN weight_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 293.745000 437.430000 293.885000 437.570000 ;
    END
  END weight_i[2]
  PIN weight_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 294.585000 437.430000 294.725000 437.570000 ;
    END
  END weight_i[1]
  PIN weight_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 295.425000 437.430000 295.565000 437.570000 ;
    END
  END weight_i[0]
  PIN dout_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 264.315000 368.980000 264.455000 ;
    END
  END dout_o[159]
  PIN dout_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 263.745000 368.980000 263.885000 ;
    END
  END dout_o[158]
  PIN dout_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 263.175000 368.980000 263.315000 ;
    END
  END dout_o[157]
  PIN dout_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 262.605000 368.980000 262.745000 ;
    END
  END dout_o[156]
  PIN dout_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 262.035000 368.980000 262.175000 ;
    END
  END dout_o[155]
  PIN dout_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 261.465000 368.980000 261.605000 ;
    END
  END dout_o[154]
  PIN dout_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 260.895000 368.980000 261.035000 ;
    END
  END dout_o[153]
  PIN dout_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 260.325000 368.980000 260.465000 ;
    END
  END dout_o[152]
  PIN dout_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 259.755000 368.980000 259.895000 ;
    END
  END dout_o[151]
  PIN dout_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 259.185000 368.980000 259.325000 ;
    END
  END dout_o[150]
  PIN dout_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 258.615000 368.980000 258.755000 ;
    END
  END dout_o[149]
  PIN dout_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 258.045000 368.980000 258.185000 ;
    END
  END dout_o[148]
  PIN dout_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 257.475000 368.980000 257.615000 ;
    END
  END dout_o[147]
  PIN dout_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 256.905000 368.980000 257.045000 ;
    END
  END dout_o[146]
  PIN dout_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 256.335000 368.980000 256.475000 ;
    END
  END dout_o[145]
  PIN dout_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 255.765000 368.980000 255.905000 ;
    END
  END dout_o[144]
  PIN dout_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 255.195000 368.980000 255.335000 ;
    END
  END dout_o[143]
  PIN dout_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 254.625000 368.980000 254.765000 ;
    END
  END dout_o[142]
  PIN dout_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 254.055000 368.980000 254.195000 ;
    END
  END dout_o[141]
  PIN dout_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 253.485000 368.980000 253.625000 ;
    END
  END dout_o[140]
  PIN dout_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 252.915000 368.980000 253.055000 ;
    END
  END dout_o[139]
  PIN dout_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 252.345000 368.980000 252.485000 ;
    END
  END dout_o[138]
  PIN dout_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 251.775000 368.980000 251.915000 ;
    END
  END dout_o[137]
  PIN dout_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 251.205000 368.980000 251.345000 ;
    END
  END dout_o[136]
  PIN dout_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 250.635000 368.980000 250.775000 ;
    END
  END dout_o[135]
  PIN dout_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 250.065000 368.980000 250.205000 ;
    END
  END dout_o[134]
  PIN dout_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 249.495000 368.980000 249.635000 ;
    END
  END dout_o[133]
  PIN dout_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 248.925000 368.980000 249.065000 ;
    END
  END dout_o[132]
  PIN dout_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 248.355000 368.980000 248.495000 ;
    END
  END dout_o[131]
  PIN dout_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 247.785000 368.980000 247.925000 ;
    END
  END dout_o[130]
  PIN dout_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 247.215000 368.980000 247.355000 ;
    END
  END dout_o[129]
  PIN dout_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 246.645000 368.980000 246.785000 ;
    END
  END dout_o[128]
  PIN dout_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 246.075000 368.980000 246.215000 ;
    END
  END dout_o[127]
  PIN dout_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 245.505000 368.980000 245.645000 ;
    END
  END dout_o[126]
  PIN dout_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 244.935000 368.980000 245.075000 ;
    END
  END dout_o[125]
  PIN dout_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 244.365000 368.980000 244.505000 ;
    END
  END dout_o[124]
  PIN dout_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 243.795000 368.980000 243.935000 ;
    END
  END dout_o[123]
  PIN dout_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 243.225000 368.980000 243.365000 ;
    END
  END dout_o[122]
  PIN dout_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 242.655000 368.980000 242.795000 ;
    END
  END dout_o[121]
  PIN dout_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 242.085000 368.980000 242.225000 ;
    END
  END dout_o[120]
  PIN dout_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 241.515000 368.980000 241.655000 ;
    END
  END dout_o[119]
  PIN dout_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 240.945000 368.980000 241.085000 ;
    END
  END dout_o[118]
  PIN dout_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 240.375000 368.980000 240.515000 ;
    END
  END dout_o[117]
  PIN dout_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 239.805000 368.980000 239.945000 ;
    END
  END dout_o[116]
  PIN dout_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 239.235000 368.980000 239.375000 ;
    END
  END dout_o[115]
  PIN dout_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 238.665000 368.980000 238.805000 ;
    END
  END dout_o[114]
  PIN dout_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 238.095000 368.980000 238.235000 ;
    END
  END dout_o[113]
  PIN dout_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 237.525000 368.980000 237.665000 ;
    END
  END dout_o[112]
  PIN dout_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 236.955000 368.980000 237.095000 ;
    END
  END dout_o[111]
  PIN dout_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 236.385000 368.980000 236.525000 ;
    END
  END dout_o[110]
  PIN dout_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 235.815000 368.980000 235.955000 ;
    END
  END dout_o[109]
  PIN dout_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 235.245000 368.980000 235.385000 ;
    END
  END dout_o[108]
  PIN dout_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 234.675000 368.980000 234.815000 ;
    END
  END dout_o[107]
  PIN dout_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 234.105000 368.980000 234.245000 ;
    END
  END dout_o[106]
  PIN dout_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 233.535000 368.980000 233.675000 ;
    END
  END dout_o[105]
  PIN dout_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 232.965000 368.980000 233.105000 ;
    END
  END dout_o[104]
  PIN dout_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 232.395000 368.980000 232.535000 ;
    END
  END dout_o[103]
  PIN dout_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 231.825000 368.980000 231.965000 ;
    END
  END dout_o[102]
  PIN dout_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 231.255000 368.980000 231.395000 ;
    END
  END dout_o[101]
  PIN dout_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 230.685000 368.980000 230.825000 ;
    END
  END dout_o[100]
  PIN dout_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 230.115000 368.980000 230.255000 ;
    END
  END dout_o[99]
  PIN dout_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 229.545000 368.980000 229.685000 ;
    END
  END dout_o[98]
  PIN dout_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 228.975000 368.980000 229.115000 ;
    END
  END dout_o[97]
  PIN dout_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 228.405000 368.980000 228.545000 ;
    END
  END dout_o[96]
  PIN dout_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 227.835000 368.980000 227.975000 ;
    END
  END dout_o[95]
  PIN dout_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 227.265000 368.980000 227.405000 ;
    END
  END dout_o[94]
  PIN dout_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 226.695000 368.980000 226.835000 ;
    END
  END dout_o[93]
  PIN dout_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 226.125000 368.980000 226.265000 ;
    END
  END dout_o[92]
  PIN dout_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 225.555000 368.980000 225.695000 ;
    END
  END dout_o[91]
  PIN dout_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 224.985000 368.980000 225.125000 ;
    END
  END dout_o[90]
  PIN dout_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 224.415000 368.980000 224.555000 ;
    END
  END dout_o[89]
  PIN dout_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 223.845000 368.980000 223.985000 ;
    END
  END dout_o[88]
  PIN dout_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 223.275000 368.980000 223.415000 ;
    END
  END dout_o[87]
  PIN dout_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 222.705000 368.980000 222.845000 ;
    END
  END dout_o[86]
  PIN dout_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 222.135000 368.980000 222.275000 ;
    END
  END dout_o[85]
  PIN dout_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 221.565000 368.980000 221.705000 ;
    END
  END dout_o[84]
  PIN dout_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 220.995000 368.980000 221.135000 ;
    END
  END dout_o[83]
  PIN dout_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 220.425000 368.980000 220.565000 ;
    END
  END dout_o[82]
  PIN dout_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 219.855000 368.980000 219.995000 ;
    END
  END dout_o[81]
  PIN dout_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 219.285000 368.980000 219.425000 ;
    END
  END dout_o[80]
  PIN dout_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 218.715000 368.980000 218.855000 ;
    END
  END dout_o[79]
  PIN dout_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 218.145000 368.980000 218.285000 ;
    END
  END dout_o[78]
  PIN dout_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 217.575000 368.980000 217.715000 ;
    END
  END dout_o[77]
  PIN dout_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 217.005000 368.980000 217.145000 ;
    END
  END dout_o[76]
  PIN dout_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 216.435000 368.980000 216.575000 ;
    END
  END dout_o[75]
  PIN dout_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 215.865000 368.980000 216.005000 ;
    END
  END dout_o[74]
  PIN dout_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 215.295000 368.980000 215.435000 ;
    END
  END dout_o[73]
  PIN dout_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 214.725000 368.980000 214.865000 ;
    END
  END dout_o[72]
  PIN dout_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 214.155000 368.980000 214.295000 ;
    END
  END dout_o[71]
  PIN dout_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 213.585000 368.980000 213.725000 ;
    END
  END dout_o[70]
  PIN dout_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 213.015000 368.980000 213.155000 ;
    END
  END dout_o[69]
  PIN dout_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 212.445000 368.980000 212.585000 ;
    END
  END dout_o[68]
  PIN dout_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 211.875000 368.980000 212.015000 ;
    END
  END dout_o[67]
  PIN dout_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 211.305000 368.980000 211.445000 ;
    END
  END dout_o[66]
  PIN dout_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 210.735000 368.980000 210.875000 ;
    END
  END dout_o[65]
  PIN dout_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 210.165000 368.980000 210.305000 ;
    END
  END dout_o[64]
  PIN dout_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 209.595000 368.980000 209.735000 ;
    END
  END dout_o[63]
  PIN dout_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 209.025000 368.980000 209.165000 ;
    END
  END dout_o[62]
  PIN dout_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 208.455000 368.980000 208.595000 ;
    END
  END dout_o[61]
  PIN dout_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 207.885000 368.980000 208.025000 ;
    END
  END dout_o[60]
  PIN dout_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 207.315000 368.980000 207.455000 ;
    END
  END dout_o[59]
  PIN dout_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 206.745000 368.980000 206.885000 ;
    END
  END dout_o[58]
  PIN dout_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 206.175000 368.980000 206.315000 ;
    END
  END dout_o[57]
  PIN dout_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 205.605000 368.980000 205.745000 ;
    END
  END dout_o[56]
  PIN dout_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 205.035000 368.980000 205.175000 ;
    END
  END dout_o[55]
  PIN dout_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 204.465000 368.980000 204.605000 ;
    END
  END dout_o[54]
  PIN dout_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 203.895000 368.980000 204.035000 ;
    END
  END dout_o[53]
  PIN dout_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 203.325000 368.980000 203.465000 ;
    END
  END dout_o[52]
  PIN dout_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 202.755000 368.980000 202.895000 ;
    END
  END dout_o[51]
  PIN dout_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 202.185000 368.980000 202.325000 ;
    END
  END dout_o[50]
  PIN dout_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 201.615000 368.980000 201.755000 ;
    END
  END dout_o[49]
  PIN dout_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 201.045000 368.980000 201.185000 ;
    END
  END dout_o[48]
  PIN dout_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 200.475000 368.980000 200.615000 ;
    END
  END dout_o[47]
  PIN dout_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 199.905000 368.980000 200.045000 ;
    END
  END dout_o[46]
  PIN dout_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 199.335000 368.980000 199.475000 ;
    END
  END dout_o[45]
  PIN dout_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 198.765000 368.980000 198.905000 ;
    END
  END dout_o[44]
  PIN dout_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 198.195000 368.980000 198.335000 ;
    END
  END dout_o[43]
  PIN dout_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 197.625000 368.980000 197.765000 ;
    END
  END dout_o[42]
  PIN dout_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 197.055000 368.980000 197.195000 ;
    END
  END dout_o[41]
  PIN dout_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 196.485000 368.980000 196.625000 ;
    END
  END dout_o[40]
  PIN dout_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 195.915000 368.980000 196.055000 ;
    END
  END dout_o[39]
  PIN dout_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 195.345000 368.980000 195.485000 ;
    END
  END dout_o[38]
  PIN dout_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 194.775000 368.980000 194.915000 ;
    END
  END dout_o[37]
  PIN dout_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 194.205000 368.980000 194.345000 ;
    END
  END dout_o[36]
  PIN dout_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 193.635000 368.980000 193.775000 ;
    END
  END dout_o[35]
  PIN dout_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 193.065000 368.980000 193.205000 ;
    END
  END dout_o[34]
  PIN dout_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 192.495000 368.980000 192.635000 ;
    END
  END dout_o[33]
  PIN dout_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 191.925000 368.980000 192.065000 ;
    END
  END dout_o[32]
  PIN dout_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 191.355000 368.980000 191.495000 ;
    END
  END dout_o[31]
  PIN dout_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 190.785000 368.980000 190.925000 ;
    END
  END dout_o[30]
  PIN dout_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 190.215000 368.980000 190.355000 ;
    END
  END dout_o[29]
  PIN dout_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 189.645000 368.980000 189.785000 ;
    END
  END dout_o[28]
  PIN dout_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 189.075000 368.980000 189.215000 ;
    END
  END dout_o[27]
  PIN dout_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 188.505000 368.980000 188.645000 ;
    END
  END dout_o[26]
  PIN dout_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 187.935000 368.980000 188.075000 ;
    END
  END dout_o[25]
  PIN dout_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 187.365000 368.980000 187.505000 ;
    END
  END dout_o[24]
  PIN dout_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 186.795000 368.980000 186.935000 ;
    END
  END dout_o[23]
  PIN dout_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 186.225000 368.980000 186.365000 ;
    END
  END dout_o[22]
  PIN dout_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 185.655000 368.980000 185.795000 ;
    END
  END dout_o[21]
  PIN dout_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 185.085000 368.980000 185.225000 ;
    END
  END dout_o[20]
  PIN dout_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 184.515000 368.980000 184.655000 ;
    END
  END dout_o[19]
  PIN dout_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 183.945000 368.980000 184.085000 ;
    END
  END dout_o[18]
  PIN dout_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 183.375000 368.980000 183.515000 ;
    END
  END dout_o[17]
  PIN dout_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 182.805000 368.980000 182.945000 ;
    END
  END dout_o[16]
  PIN dout_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 182.235000 368.980000 182.375000 ;
    END
  END dout_o[15]
  PIN dout_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 181.665000 368.980000 181.805000 ;
    END
  END dout_o[14]
  PIN dout_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 181.095000 368.980000 181.235000 ;
    END
  END dout_o[13]
  PIN dout_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 180.525000 368.980000 180.665000 ;
    END
  END dout_o[12]
  PIN dout_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 179.955000 368.980000 180.095000 ;
    END
  END dout_o[11]
  PIN dout_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 179.385000 368.980000 179.525000 ;
    END
  END dout_o[10]
  PIN dout_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 178.815000 368.980000 178.955000 ;
    END
  END dout_o[9]
  PIN dout_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 178.245000 368.980000 178.385000 ;
    END
  END dout_o[8]
  PIN dout_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 177.675000 368.980000 177.815000 ;
    END
  END dout_o[7]
  PIN dout_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 177.105000 368.980000 177.245000 ;
    END
  END dout_o[6]
  PIN dout_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 176.535000 368.980000 176.675000 ;
    END
  END dout_o[5]
  PIN dout_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 175.965000 368.980000 176.105000 ;
    END
  END dout_o[4]
  PIN dout_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 175.395000 368.980000 175.535000 ;
    END
  END dout_o[3]
  PIN dout_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 174.825000 368.980000 174.965000 ;
    END
  END dout_o[2]
  PIN dout_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 174.255000 368.980000 174.395000 ;
    END
  END dout_o[1]
  PIN dout_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 368.840000 173.685000 368.980000 173.825000 ;
    END
  END dout_o[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal4 ;
      RECT 295.705000 437.290000 368.980000 437.570000 ;
      RECT 294.865000 437.290000 295.285000 437.570000 ;
      RECT 294.025000 437.290000 294.445000 437.570000 ;
      RECT 293.185000 437.290000 293.605000 437.570000 ;
      RECT 292.345000 437.290000 292.765000 437.570000 ;
      RECT 291.505000 437.290000 291.925000 437.570000 ;
      RECT 290.665000 437.290000 291.085000 437.570000 ;
      RECT 289.825000 437.290000 290.245000 437.570000 ;
      RECT 288.985000 437.290000 289.405000 437.570000 ;
      RECT 288.145000 437.290000 288.565000 437.570000 ;
      RECT 287.305000 437.290000 287.725000 437.570000 ;
      RECT 286.465000 437.290000 286.885000 437.570000 ;
      RECT 285.625000 437.290000 286.045000 437.570000 ;
      RECT 284.785000 437.290000 285.205000 437.570000 ;
      RECT 283.945000 437.290000 284.365000 437.570000 ;
      RECT 283.105000 437.290000 283.525000 437.570000 ;
      RECT 282.265000 437.290000 282.685000 437.570000 ;
      RECT 281.425000 437.290000 281.845000 437.570000 ;
      RECT 280.585000 437.290000 281.005000 437.570000 ;
      RECT 279.745000 437.290000 280.165000 437.570000 ;
      RECT 278.905000 437.290000 279.325000 437.570000 ;
      RECT 278.065000 437.290000 278.485000 437.570000 ;
      RECT 277.225000 437.290000 277.645000 437.570000 ;
      RECT 276.385000 437.290000 276.805000 437.570000 ;
      RECT 275.545000 437.290000 275.965000 437.570000 ;
      RECT 274.705000 437.290000 275.125000 437.570000 ;
      RECT 273.865000 437.290000 274.285000 437.570000 ;
      RECT 273.025000 437.290000 273.445000 437.570000 ;
      RECT 272.185000 437.290000 272.605000 437.570000 ;
      RECT 271.345000 437.290000 271.765000 437.570000 ;
      RECT 270.505000 437.290000 270.925000 437.570000 ;
      RECT 269.665000 437.290000 270.085000 437.570000 ;
      RECT 268.825000 437.290000 269.245000 437.570000 ;
      RECT 267.985000 437.290000 268.405000 437.570000 ;
      RECT 267.145000 437.290000 267.565000 437.570000 ;
      RECT 266.305000 437.290000 266.725000 437.570000 ;
      RECT 265.465000 437.290000 265.885000 437.570000 ;
      RECT 264.625000 437.290000 265.045000 437.570000 ;
      RECT 263.785000 437.290000 264.205000 437.570000 ;
      RECT 262.945000 437.290000 263.365000 437.570000 ;
      RECT 262.105000 437.290000 262.525000 437.570000 ;
      RECT 261.265000 437.290000 261.685000 437.570000 ;
      RECT 260.425000 437.290000 260.845000 437.570000 ;
      RECT 259.585000 437.290000 260.005000 437.570000 ;
      RECT 258.745000 437.290000 259.165000 437.570000 ;
      RECT 257.905000 437.290000 258.325000 437.570000 ;
      RECT 257.065000 437.290000 257.485000 437.570000 ;
      RECT 256.225000 437.290000 256.645000 437.570000 ;
      RECT 255.385000 437.290000 255.805000 437.570000 ;
      RECT 254.545000 437.290000 254.965000 437.570000 ;
      RECT 253.705000 437.290000 254.125000 437.570000 ;
      RECT 252.865000 437.290000 253.285000 437.570000 ;
      RECT 252.025000 437.290000 252.445000 437.570000 ;
      RECT 251.185000 437.290000 251.605000 437.570000 ;
      RECT 250.345000 437.290000 250.765000 437.570000 ;
      RECT 249.505000 437.290000 249.925000 437.570000 ;
      RECT 248.665000 437.290000 249.085000 437.570000 ;
      RECT 247.825000 437.290000 248.245000 437.570000 ;
      RECT 246.985000 437.290000 247.405000 437.570000 ;
      RECT 246.145000 437.290000 246.565000 437.570000 ;
      RECT 245.305000 437.290000 245.725000 437.570000 ;
      RECT 244.465000 437.290000 244.885000 437.570000 ;
      RECT 243.625000 437.290000 244.045000 437.570000 ;
      RECT 242.785000 437.290000 243.205000 437.570000 ;
      RECT 241.945000 437.290000 242.365000 437.570000 ;
      RECT 241.105000 437.290000 241.525000 437.570000 ;
      RECT 240.265000 437.290000 240.685000 437.570000 ;
      RECT 239.425000 437.290000 239.845000 437.570000 ;
      RECT 238.585000 437.290000 239.005000 437.570000 ;
      RECT 237.745000 437.290000 238.165000 437.570000 ;
      RECT 236.905000 437.290000 237.325000 437.570000 ;
      RECT 236.065000 437.290000 236.485000 437.570000 ;
      RECT 235.225000 437.290000 235.645000 437.570000 ;
      RECT 234.385000 437.290000 234.805000 437.570000 ;
      RECT 233.545000 437.290000 233.965000 437.570000 ;
      RECT 232.705000 437.290000 233.125000 437.570000 ;
      RECT 231.865000 437.290000 232.285000 437.570000 ;
      RECT 231.025000 437.290000 231.445000 437.570000 ;
      RECT 230.185000 437.290000 230.605000 437.570000 ;
      RECT 229.345000 437.290000 229.765000 437.570000 ;
      RECT 228.505000 437.290000 228.925000 437.570000 ;
      RECT 227.665000 437.290000 228.085000 437.570000 ;
      RECT 226.825000 437.290000 227.245000 437.570000 ;
      RECT 225.985000 437.290000 226.405000 437.570000 ;
      RECT 225.145000 437.290000 225.565000 437.570000 ;
      RECT 224.305000 437.290000 224.725000 437.570000 ;
      RECT 223.465000 437.290000 223.885000 437.570000 ;
      RECT 222.625000 437.290000 223.045000 437.570000 ;
      RECT 221.785000 437.290000 222.205000 437.570000 ;
      RECT 220.945000 437.290000 221.365000 437.570000 ;
      RECT 220.105000 437.290000 220.525000 437.570000 ;
      RECT 219.265000 437.290000 219.685000 437.570000 ;
      RECT 218.425000 437.290000 218.845000 437.570000 ;
      RECT 217.585000 437.290000 218.005000 437.570000 ;
      RECT 216.745000 437.290000 217.165000 437.570000 ;
      RECT 215.905000 437.290000 216.325000 437.570000 ;
      RECT 215.065000 437.290000 215.485000 437.570000 ;
      RECT 214.225000 437.290000 214.645000 437.570000 ;
      RECT 213.385000 437.290000 213.805000 437.570000 ;
      RECT 212.545000 437.290000 212.965000 437.570000 ;
      RECT 211.705000 437.290000 212.125000 437.570000 ;
      RECT 210.865000 437.290000 211.285000 437.570000 ;
      RECT 210.025000 437.290000 210.445000 437.570000 ;
      RECT 209.185000 437.290000 209.605000 437.570000 ;
      RECT 208.345000 437.290000 208.765000 437.570000 ;
      RECT 207.505000 437.290000 207.925000 437.570000 ;
      RECT 206.665000 437.290000 207.085000 437.570000 ;
      RECT 205.825000 437.290000 206.245000 437.570000 ;
      RECT 204.985000 437.290000 205.405000 437.570000 ;
      RECT 204.145000 437.290000 204.565000 437.570000 ;
      RECT 203.305000 437.290000 203.725000 437.570000 ;
      RECT 202.465000 437.290000 202.885000 437.570000 ;
      RECT 201.625000 437.290000 202.045000 437.570000 ;
      RECT 200.785000 437.290000 201.205000 437.570000 ;
      RECT 199.945000 437.290000 200.365000 437.570000 ;
      RECT 199.105000 437.290000 199.525000 437.570000 ;
      RECT 198.265000 437.290000 198.685000 437.570000 ;
      RECT 197.425000 437.290000 197.845000 437.570000 ;
      RECT 196.585000 437.290000 197.005000 437.570000 ;
      RECT 195.745000 437.290000 196.165000 437.570000 ;
      RECT 194.905000 437.290000 195.325000 437.570000 ;
      RECT 194.065000 437.290000 194.485000 437.570000 ;
      RECT 193.225000 437.290000 193.645000 437.570000 ;
      RECT 192.385000 437.290000 192.805000 437.570000 ;
      RECT 191.545000 437.290000 191.965000 437.570000 ;
      RECT 190.705000 437.290000 191.125000 437.570000 ;
      RECT 189.865000 437.290000 190.285000 437.570000 ;
      RECT 189.025000 437.290000 189.445000 437.570000 ;
      RECT 188.185000 437.290000 188.605000 437.570000 ;
      RECT 187.345000 437.290000 187.765000 437.570000 ;
      RECT 186.505000 437.290000 186.925000 437.570000 ;
      RECT 185.665000 437.290000 186.085000 437.570000 ;
      RECT 184.825000 437.290000 185.245000 437.570000 ;
      RECT 183.985000 437.290000 184.405000 437.570000 ;
      RECT 183.145000 437.290000 183.565000 437.570000 ;
      RECT 182.305000 437.290000 182.725000 437.570000 ;
      RECT 181.465000 437.290000 181.885000 437.570000 ;
      RECT 180.625000 437.290000 181.045000 437.570000 ;
      RECT 179.785000 437.290000 180.205000 437.570000 ;
      RECT 178.945000 437.290000 179.365000 437.570000 ;
      RECT 178.105000 437.290000 178.525000 437.570000 ;
      RECT 177.265000 437.290000 177.685000 437.570000 ;
      RECT 176.425000 437.290000 176.845000 437.570000 ;
      RECT 175.585000 437.290000 176.005000 437.570000 ;
      RECT 174.745000 437.290000 175.165000 437.570000 ;
      RECT 173.905000 437.290000 174.325000 437.570000 ;
      RECT 173.065000 437.290000 173.485000 437.570000 ;
      RECT 172.225000 437.290000 172.645000 437.570000 ;
      RECT 171.385000 437.290000 171.805000 437.570000 ;
      RECT 170.545000 437.290000 170.965000 437.570000 ;
      RECT 169.705000 437.290000 170.125000 437.570000 ;
      RECT 168.865000 437.290000 169.285000 437.570000 ;
      RECT 168.025000 437.290000 168.445000 437.570000 ;
      RECT 167.185000 437.290000 167.605000 437.570000 ;
      RECT 166.345000 437.290000 166.765000 437.570000 ;
      RECT 165.505000 437.290000 165.925000 437.570000 ;
      RECT 164.665000 437.290000 165.085000 437.570000 ;
      RECT 163.825000 437.290000 164.245000 437.570000 ;
      RECT 162.985000 437.290000 163.405000 437.570000 ;
      RECT 162.145000 437.290000 162.565000 437.570000 ;
      RECT 161.305000 437.290000 161.725000 437.570000 ;
      RECT 160.465000 437.290000 160.885000 437.570000 ;
      RECT 159.625000 437.290000 160.045000 437.570000 ;
      RECT 158.785000 437.290000 159.205000 437.570000 ;
      RECT 157.945000 437.290000 158.365000 437.570000 ;
      RECT 157.105000 437.290000 157.525000 437.570000 ;
      RECT 156.265000 437.290000 156.685000 437.570000 ;
      RECT 155.425000 437.290000 155.845000 437.570000 ;
      RECT 154.585000 437.290000 155.005000 437.570000 ;
      RECT 153.745000 437.290000 154.165000 437.570000 ;
      RECT 152.905000 437.290000 153.325000 437.570000 ;
      RECT 152.065000 437.290000 152.485000 437.570000 ;
      RECT 151.225000 437.290000 151.645000 437.570000 ;
      RECT 150.385000 437.290000 150.805000 437.570000 ;
      RECT 149.545000 437.290000 149.965000 437.570000 ;
      RECT 148.705000 437.290000 149.125000 437.570000 ;
      RECT 147.865000 437.290000 148.285000 437.570000 ;
      RECT 147.025000 437.290000 147.445000 437.570000 ;
      RECT 146.185000 437.290000 146.605000 437.570000 ;
      RECT 145.345000 437.290000 145.765000 437.570000 ;
      RECT 144.505000 437.290000 144.925000 437.570000 ;
      RECT 143.665000 437.290000 144.085000 437.570000 ;
      RECT 142.825000 437.290000 143.245000 437.570000 ;
      RECT 141.985000 437.290000 142.405000 437.570000 ;
      RECT 141.145000 437.290000 141.565000 437.570000 ;
      RECT 140.305000 437.290000 140.725000 437.570000 ;
      RECT 139.465000 437.290000 139.885000 437.570000 ;
      RECT 138.625000 437.290000 139.045000 437.570000 ;
      RECT 137.785000 437.290000 138.205000 437.570000 ;
      RECT 136.945000 437.290000 137.365000 437.570000 ;
      RECT 136.105000 437.290000 136.525000 437.570000 ;
      RECT 135.265000 437.290000 135.685000 437.570000 ;
      RECT 134.425000 437.290000 134.845000 437.570000 ;
      RECT 133.585000 437.290000 134.005000 437.570000 ;
      RECT 132.745000 437.290000 133.165000 437.570000 ;
      RECT 131.905000 437.290000 132.325000 437.570000 ;
      RECT 131.065000 437.290000 131.485000 437.570000 ;
      RECT 130.225000 437.290000 130.645000 437.570000 ;
      RECT 129.385000 437.290000 129.805000 437.570000 ;
      RECT 128.545000 437.290000 128.965000 437.570000 ;
      RECT 127.705000 437.290000 128.125000 437.570000 ;
      RECT 126.865000 437.290000 127.285000 437.570000 ;
      RECT 126.025000 437.290000 126.445000 437.570000 ;
      RECT 125.185000 437.290000 125.605000 437.570000 ;
      RECT 124.345000 437.290000 124.765000 437.570000 ;
      RECT 123.505000 437.290000 123.925000 437.570000 ;
      RECT 122.665000 437.290000 123.085000 437.570000 ;
      RECT 121.825000 437.290000 122.245000 437.570000 ;
      RECT 120.985000 437.290000 121.405000 437.570000 ;
      RECT 120.145000 437.290000 120.565000 437.570000 ;
      RECT 119.305000 437.290000 119.725000 437.570000 ;
      RECT 118.465000 437.290000 118.885000 437.570000 ;
      RECT 117.625000 437.290000 118.045000 437.570000 ;
      RECT 116.785000 437.290000 117.205000 437.570000 ;
      RECT 115.945000 437.290000 116.365000 437.570000 ;
      RECT 115.105000 437.290000 115.525000 437.570000 ;
      RECT 114.265000 437.290000 114.685000 437.570000 ;
      RECT 113.425000 437.290000 113.845000 437.570000 ;
      RECT 112.585000 437.290000 113.005000 437.570000 ;
      RECT 111.745000 437.290000 112.165000 437.570000 ;
      RECT 110.905000 437.290000 111.325000 437.570000 ;
      RECT 110.065000 437.290000 110.485000 437.570000 ;
      RECT 109.225000 437.290000 109.645000 437.570000 ;
      RECT 108.385000 437.290000 108.805000 437.570000 ;
      RECT 107.545000 437.290000 107.965000 437.570000 ;
      RECT 106.705000 437.290000 107.125000 437.570000 ;
      RECT 105.865000 437.290000 106.285000 437.570000 ;
      RECT 105.025000 437.290000 105.445000 437.570000 ;
      RECT 104.185000 437.290000 104.605000 437.570000 ;
      RECT 103.345000 437.290000 103.765000 437.570000 ;
      RECT 102.505000 437.290000 102.925000 437.570000 ;
      RECT 101.665000 437.290000 102.085000 437.570000 ;
      RECT 100.825000 437.290000 101.245000 437.570000 ;
      RECT 99.985000 437.290000 100.405000 437.570000 ;
      RECT 99.145000 437.290000 99.565000 437.570000 ;
      RECT 98.305000 437.290000 98.725000 437.570000 ;
      RECT 97.465000 437.290000 97.885000 437.570000 ;
      RECT 96.625000 437.290000 97.045000 437.570000 ;
      RECT 95.785000 437.290000 96.205000 437.570000 ;
      RECT 94.945000 437.290000 95.365000 437.570000 ;
      RECT 94.105000 437.290000 94.525000 437.570000 ;
      RECT 93.265000 437.290000 93.685000 437.570000 ;
      RECT 92.425000 437.290000 92.845000 437.570000 ;
      RECT 91.585000 437.290000 92.005000 437.570000 ;
      RECT 90.745000 437.290000 91.165000 437.570000 ;
      RECT 89.905000 437.290000 90.325000 437.570000 ;
      RECT 89.065000 437.290000 89.485000 437.570000 ;
      RECT 88.225000 437.290000 88.645000 437.570000 ;
      RECT 87.385000 437.290000 87.805000 437.570000 ;
      RECT 86.545000 437.290000 86.965000 437.570000 ;
      RECT 85.705000 437.290000 86.125000 437.570000 ;
      RECT 84.865000 437.290000 85.285000 437.570000 ;
      RECT 84.025000 437.290000 84.445000 437.570000 ;
      RECT 83.185000 437.290000 83.605000 437.570000 ;
      RECT 82.345000 437.290000 82.765000 437.570000 ;
      RECT 81.505000 437.290000 81.925000 437.570000 ;
      RECT 80.665000 437.290000 81.085000 437.570000 ;
      RECT 79.825000 437.290000 80.245000 437.570000 ;
      RECT 78.985000 437.290000 79.405000 437.570000 ;
      RECT 78.145000 437.290000 78.565000 437.570000 ;
      RECT 77.305000 437.290000 77.725000 437.570000 ;
      RECT 76.465000 437.290000 76.885000 437.570000 ;
      RECT 75.625000 437.290000 76.045000 437.570000 ;
      RECT 74.785000 437.290000 75.205000 437.570000 ;
      RECT 73.945000 437.290000 74.365000 437.570000 ;
      RECT 73.105000 437.290000 73.525000 437.570000 ;
      RECT 0.000000 437.290000 72.685000 437.570000 ;
      RECT 0.000000 292.905000 368.980000 437.290000 ;
      RECT 0.280000 292.485000 368.980000 292.905000 ;
      RECT 0.000000 292.335000 368.980000 292.485000 ;
      RECT 0.280000 291.915000 368.980000 292.335000 ;
      RECT 0.000000 291.765000 368.980000 291.915000 ;
      RECT 0.280000 291.345000 368.980000 291.765000 ;
      RECT 0.000000 291.195000 368.980000 291.345000 ;
      RECT 0.280000 290.775000 368.980000 291.195000 ;
      RECT 0.000000 290.625000 368.980000 290.775000 ;
      RECT 0.280000 290.205000 368.980000 290.625000 ;
      RECT 0.000000 290.055000 368.980000 290.205000 ;
      RECT 0.280000 289.635000 368.980000 290.055000 ;
      RECT 0.000000 289.485000 368.980000 289.635000 ;
      RECT 0.280000 289.065000 368.980000 289.485000 ;
      RECT 0.000000 288.915000 368.980000 289.065000 ;
      RECT 0.280000 288.495000 368.980000 288.915000 ;
      RECT 0.000000 288.345000 368.980000 288.495000 ;
      RECT 0.280000 287.925000 368.980000 288.345000 ;
      RECT 0.000000 287.775000 368.980000 287.925000 ;
      RECT 0.280000 287.355000 368.980000 287.775000 ;
      RECT 0.000000 287.205000 368.980000 287.355000 ;
      RECT 0.280000 286.785000 368.980000 287.205000 ;
      RECT 0.000000 286.635000 368.980000 286.785000 ;
      RECT 0.280000 286.215000 368.980000 286.635000 ;
      RECT 0.000000 286.065000 368.980000 286.215000 ;
      RECT 0.280000 285.645000 368.980000 286.065000 ;
      RECT 0.000000 285.495000 368.980000 285.645000 ;
      RECT 0.280000 285.075000 368.980000 285.495000 ;
      RECT 0.000000 284.925000 368.980000 285.075000 ;
      RECT 0.280000 284.505000 368.980000 284.925000 ;
      RECT 0.000000 284.355000 368.980000 284.505000 ;
      RECT 0.280000 283.935000 368.980000 284.355000 ;
      RECT 0.000000 283.785000 368.980000 283.935000 ;
      RECT 0.280000 283.365000 368.980000 283.785000 ;
      RECT 0.000000 283.215000 368.980000 283.365000 ;
      RECT 0.280000 282.795000 368.980000 283.215000 ;
      RECT 0.000000 282.645000 368.980000 282.795000 ;
      RECT 0.280000 282.225000 368.980000 282.645000 ;
      RECT 0.000000 282.075000 368.980000 282.225000 ;
      RECT 0.280000 281.655000 368.980000 282.075000 ;
      RECT 0.000000 281.505000 368.980000 281.655000 ;
      RECT 0.280000 281.085000 368.980000 281.505000 ;
      RECT 0.000000 280.935000 368.980000 281.085000 ;
      RECT 0.280000 280.515000 368.980000 280.935000 ;
      RECT 0.000000 280.365000 368.980000 280.515000 ;
      RECT 0.280000 279.945000 368.980000 280.365000 ;
      RECT 0.000000 279.795000 368.980000 279.945000 ;
      RECT 0.280000 279.375000 368.980000 279.795000 ;
      RECT 0.000000 279.225000 368.980000 279.375000 ;
      RECT 0.280000 278.805000 368.980000 279.225000 ;
      RECT 0.000000 278.655000 368.980000 278.805000 ;
      RECT 0.280000 278.235000 368.980000 278.655000 ;
      RECT 0.000000 278.085000 368.980000 278.235000 ;
      RECT 0.280000 277.665000 368.980000 278.085000 ;
      RECT 0.000000 277.515000 368.980000 277.665000 ;
      RECT 0.280000 277.095000 368.980000 277.515000 ;
      RECT 0.000000 276.945000 368.980000 277.095000 ;
      RECT 0.280000 276.525000 368.980000 276.945000 ;
      RECT 0.000000 276.375000 368.980000 276.525000 ;
      RECT 0.280000 275.955000 368.980000 276.375000 ;
      RECT 0.000000 275.805000 368.980000 275.955000 ;
      RECT 0.280000 275.385000 368.980000 275.805000 ;
      RECT 0.000000 275.235000 368.980000 275.385000 ;
      RECT 0.280000 274.815000 368.980000 275.235000 ;
      RECT 0.000000 274.665000 368.980000 274.815000 ;
      RECT 0.280000 274.245000 368.980000 274.665000 ;
      RECT 0.000000 274.095000 368.980000 274.245000 ;
      RECT 0.280000 273.675000 368.980000 274.095000 ;
      RECT 0.000000 273.525000 368.980000 273.675000 ;
      RECT 0.280000 273.105000 368.980000 273.525000 ;
      RECT 0.000000 272.955000 368.980000 273.105000 ;
      RECT 0.280000 272.535000 368.980000 272.955000 ;
      RECT 0.000000 272.385000 368.980000 272.535000 ;
      RECT 0.280000 271.965000 368.980000 272.385000 ;
      RECT 0.000000 271.815000 368.980000 271.965000 ;
      RECT 0.280000 271.395000 368.980000 271.815000 ;
      RECT 0.000000 271.245000 368.980000 271.395000 ;
      RECT 0.280000 270.825000 368.980000 271.245000 ;
      RECT 0.000000 270.675000 368.980000 270.825000 ;
      RECT 0.280000 270.255000 368.980000 270.675000 ;
      RECT 0.000000 270.105000 368.980000 270.255000 ;
      RECT 0.280000 269.685000 368.980000 270.105000 ;
      RECT 0.000000 269.535000 368.980000 269.685000 ;
      RECT 0.280000 269.115000 368.980000 269.535000 ;
      RECT 0.000000 268.965000 368.980000 269.115000 ;
      RECT 0.280000 268.545000 368.980000 268.965000 ;
      RECT 0.000000 268.395000 368.980000 268.545000 ;
      RECT 0.280000 267.975000 368.980000 268.395000 ;
      RECT 0.000000 267.825000 368.980000 267.975000 ;
      RECT 0.280000 267.405000 368.980000 267.825000 ;
      RECT 0.000000 267.255000 368.980000 267.405000 ;
      RECT 0.280000 266.835000 368.980000 267.255000 ;
      RECT 0.000000 266.685000 368.980000 266.835000 ;
      RECT 0.280000 266.265000 368.980000 266.685000 ;
      RECT 0.000000 266.115000 368.980000 266.265000 ;
      RECT 0.280000 265.695000 368.980000 266.115000 ;
      RECT 0.000000 265.545000 368.980000 265.695000 ;
      RECT 0.280000 265.125000 368.980000 265.545000 ;
      RECT 0.000000 264.975000 368.980000 265.125000 ;
      RECT 0.280000 264.595000 368.980000 264.975000 ;
      RECT 0.280000 264.555000 368.700000 264.595000 ;
      RECT 0.000000 264.405000 368.700000 264.555000 ;
      RECT 0.280000 264.175000 368.700000 264.405000 ;
      RECT 0.280000 264.025000 368.980000 264.175000 ;
      RECT 0.280000 263.985000 368.700000 264.025000 ;
      RECT 0.000000 263.835000 368.700000 263.985000 ;
      RECT 0.280000 263.605000 368.700000 263.835000 ;
      RECT 0.280000 263.455000 368.980000 263.605000 ;
      RECT 0.280000 263.415000 368.700000 263.455000 ;
      RECT 0.000000 263.265000 368.700000 263.415000 ;
      RECT 0.280000 263.035000 368.700000 263.265000 ;
      RECT 0.280000 262.885000 368.980000 263.035000 ;
      RECT 0.280000 262.845000 368.700000 262.885000 ;
      RECT 0.000000 262.695000 368.700000 262.845000 ;
      RECT 0.280000 262.465000 368.700000 262.695000 ;
      RECT 0.280000 262.315000 368.980000 262.465000 ;
      RECT 0.280000 262.275000 368.700000 262.315000 ;
      RECT 0.000000 262.125000 368.700000 262.275000 ;
      RECT 0.280000 261.895000 368.700000 262.125000 ;
      RECT 0.280000 261.745000 368.980000 261.895000 ;
      RECT 0.280000 261.705000 368.700000 261.745000 ;
      RECT 0.000000 261.555000 368.700000 261.705000 ;
      RECT 0.280000 261.325000 368.700000 261.555000 ;
      RECT 0.280000 261.175000 368.980000 261.325000 ;
      RECT 0.280000 261.135000 368.700000 261.175000 ;
      RECT 0.000000 260.985000 368.700000 261.135000 ;
      RECT 0.280000 260.755000 368.700000 260.985000 ;
      RECT 0.280000 260.605000 368.980000 260.755000 ;
      RECT 0.280000 260.565000 368.700000 260.605000 ;
      RECT 0.000000 260.415000 368.700000 260.565000 ;
      RECT 0.280000 260.185000 368.700000 260.415000 ;
      RECT 0.280000 260.035000 368.980000 260.185000 ;
      RECT 0.280000 259.995000 368.700000 260.035000 ;
      RECT 0.000000 259.845000 368.700000 259.995000 ;
      RECT 0.280000 259.615000 368.700000 259.845000 ;
      RECT 0.280000 259.465000 368.980000 259.615000 ;
      RECT 0.280000 259.425000 368.700000 259.465000 ;
      RECT 0.000000 259.275000 368.700000 259.425000 ;
      RECT 0.280000 259.045000 368.700000 259.275000 ;
      RECT 0.280000 258.895000 368.980000 259.045000 ;
      RECT 0.280000 258.855000 368.700000 258.895000 ;
      RECT 0.000000 258.705000 368.700000 258.855000 ;
      RECT 0.280000 258.475000 368.700000 258.705000 ;
      RECT 0.280000 258.325000 368.980000 258.475000 ;
      RECT 0.280000 258.285000 368.700000 258.325000 ;
      RECT 0.000000 258.135000 368.700000 258.285000 ;
      RECT 0.280000 257.905000 368.700000 258.135000 ;
      RECT 0.280000 257.755000 368.980000 257.905000 ;
      RECT 0.280000 257.715000 368.700000 257.755000 ;
      RECT 0.000000 257.565000 368.700000 257.715000 ;
      RECT 0.280000 257.335000 368.700000 257.565000 ;
      RECT 0.280000 257.185000 368.980000 257.335000 ;
      RECT 0.280000 257.145000 368.700000 257.185000 ;
      RECT 0.000000 256.995000 368.700000 257.145000 ;
      RECT 0.280000 256.765000 368.700000 256.995000 ;
      RECT 0.280000 256.615000 368.980000 256.765000 ;
      RECT 0.280000 256.575000 368.700000 256.615000 ;
      RECT 0.000000 256.425000 368.700000 256.575000 ;
      RECT 0.280000 256.195000 368.700000 256.425000 ;
      RECT 0.280000 256.045000 368.980000 256.195000 ;
      RECT 0.280000 256.005000 368.700000 256.045000 ;
      RECT 0.000000 255.855000 368.700000 256.005000 ;
      RECT 0.280000 255.625000 368.700000 255.855000 ;
      RECT 0.280000 255.475000 368.980000 255.625000 ;
      RECT 0.280000 255.435000 368.700000 255.475000 ;
      RECT 0.000000 255.285000 368.700000 255.435000 ;
      RECT 0.280000 255.055000 368.700000 255.285000 ;
      RECT 0.280000 254.905000 368.980000 255.055000 ;
      RECT 0.280000 254.865000 368.700000 254.905000 ;
      RECT 0.000000 254.715000 368.700000 254.865000 ;
      RECT 0.280000 254.485000 368.700000 254.715000 ;
      RECT 0.280000 254.335000 368.980000 254.485000 ;
      RECT 0.280000 254.295000 368.700000 254.335000 ;
      RECT 0.000000 254.145000 368.700000 254.295000 ;
      RECT 0.280000 253.915000 368.700000 254.145000 ;
      RECT 0.280000 253.765000 368.980000 253.915000 ;
      RECT 0.280000 253.725000 368.700000 253.765000 ;
      RECT 0.000000 253.575000 368.700000 253.725000 ;
      RECT 0.280000 253.345000 368.700000 253.575000 ;
      RECT 0.280000 253.195000 368.980000 253.345000 ;
      RECT 0.280000 253.155000 368.700000 253.195000 ;
      RECT 0.000000 253.005000 368.700000 253.155000 ;
      RECT 0.280000 252.775000 368.700000 253.005000 ;
      RECT 0.280000 252.625000 368.980000 252.775000 ;
      RECT 0.280000 252.585000 368.700000 252.625000 ;
      RECT 0.000000 252.435000 368.700000 252.585000 ;
      RECT 0.280000 252.205000 368.700000 252.435000 ;
      RECT 0.280000 252.055000 368.980000 252.205000 ;
      RECT 0.280000 252.015000 368.700000 252.055000 ;
      RECT 0.000000 251.865000 368.700000 252.015000 ;
      RECT 0.280000 251.635000 368.700000 251.865000 ;
      RECT 0.280000 251.485000 368.980000 251.635000 ;
      RECT 0.280000 251.445000 368.700000 251.485000 ;
      RECT 0.000000 251.295000 368.700000 251.445000 ;
      RECT 0.280000 251.065000 368.700000 251.295000 ;
      RECT 0.280000 250.915000 368.980000 251.065000 ;
      RECT 0.280000 250.875000 368.700000 250.915000 ;
      RECT 0.000000 250.725000 368.700000 250.875000 ;
      RECT 0.280000 250.495000 368.700000 250.725000 ;
      RECT 0.280000 250.345000 368.980000 250.495000 ;
      RECT 0.280000 250.305000 368.700000 250.345000 ;
      RECT 0.000000 250.155000 368.700000 250.305000 ;
      RECT 0.280000 249.925000 368.700000 250.155000 ;
      RECT 0.280000 249.775000 368.980000 249.925000 ;
      RECT 0.280000 249.735000 368.700000 249.775000 ;
      RECT 0.000000 249.585000 368.700000 249.735000 ;
      RECT 0.280000 249.355000 368.700000 249.585000 ;
      RECT 0.280000 249.205000 368.980000 249.355000 ;
      RECT 0.280000 249.165000 368.700000 249.205000 ;
      RECT 0.000000 249.015000 368.700000 249.165000 ;
      RECT 0.280000 248.785000 368.700000 249.015000 ;
      RECT 0.280000 248.635000 368.980000 248.785000 ;
      RECT 0.280000 248.595000 368.700000 248.635000 ;
      RECT 0.000000 248.445000 368.700000 248.595000 ;
      RECT 0.280000 248.215000 368.700000 248.445000 ;
      RECT 0.280000 248.065000 368.980000 248.215000 ;
      RECT 0.280000 248.025000 368.700000 248.065000 ;
      RECT 0.000000 247.875000 368.700000 248.025000 ;
      RECT 0.280000 247.645000 368.700000 247.875000 ;
      RECT 0.280000 247.495000 368.980000 247.645000 ;
      RECT 0.280000 247.455000 368.700000 247.495000 ;
      RECT 0.000000 247.305000 368.700000 247.455000 ;
      RECT 0.280000 247.075000 368.700000 247.305000 ;
      RECT 0.280000 246.925000 368.980000 247.075000 ;
      RECT 0.280000 246.885000 368.700000 246.925000 ;
      RECT 0.000000 246.735000 368.700000 246.885000 ;
      RECT 0.280000 246.505000 368.700000 246.735000 ;
      RECT 0.280000 246.355000 368.980000 246.505000 ;
      RECT 0.280000 246.315000 368.700000 246.355000 ;
      RECT 0.000000 246.165000 368.700000 246.315000 ;
      RECT 0.280000 245.935000 368.700000 246.165000 ;
      RECT 0.280000 245.785000 368.980000 245.935000 ;
      RECT 0.280000 245.745000 368.700000 245.785000 ;
      RECT 0.000000 245.595000 368.700000 245.745000 ;
      RECT 0.280000 245.365000 368.700000 245.595000 ;
      RECT 0.280000 245.215000 368.980000 245.365000 ;
      RECT 0.280000 245.175000 368.700000 245.215000 ;
      RECT 0.000000 245.025000 368.700000 245.175000 ;
      RECT 0.280000 244.795000 368.700000 245.025000 ;
      RECT 0.280000 244.645000 368.980000 244.795000 ;
      RECT 0.280000 244.605000 368.700000 244.645000 ;
      RECT 0.000000 244.455000 368.700000 244.605000 ;
      RECT 0.280000 244.225000 368.700000 244.455000 ;
      RECT 0.280000 244.075000 368.980000 244.225000 ;
      RECT 0.280000 244.035000 368.700000 244.075000 ;
      RECT 0.000000 243.885000 368.700000 244.035000 ;
      RECT 0.280000 243.655000 368.700000 243.885000 ;
      RECT 0.280000 243.505000 368.980000 243.655000 ;
      RECT 0.280000 243.465000 368.700000 243.505000 ;
      RECT 0.000000 243.315000 368.700000 243.465000 ;
      RECT 0.280000 243.085000 368.700000 243.315000 ;
      RECT 0.280000 242.935000 368.980000 243.085000 ;
      RECT 0.280000 242.895000 368.700000 242.935000 ;
      RECT 0.000000 242.745000 368.700000 242.895000 ;
      RECT 0.280000 242.515000 368.700000 242.745000 ;
      RECT 0.280000 242.365000 368.980000 242.515000 ;
      RECT 0.280000 242.325000 368.700000 242.365000 ;
      RECT 0.000000 242.175000 368.700000 242.325000 ;
      RECT 0.280000 241.945000 368.700000 242.175000 ;
      RECT 0.280000 241.795000 368.980000 241.945000 ;
      RECT 0.280000 241.755000 368.700000 241.795000 ;
      RECT 0.000000 241.605000 368.700000 241.755000 ;
      RECT 0.280000 241.375000 368.700000 241.605000 ;
      RECT 0.280000 241.225000 368.980000 241.375000 ;
      RECT 0.280000 241.185000 368.700000 241.225000 ;
      RECT 0.000000 241.035000 368.700000 241.185000 ;
      RECT 0.280000 240.805000 368.700000 241.035000 ;
      RECT 0.280000 240.655000 368.980000 240.805000 ;
      RECT 0.280000 240.615000 368.700000 240.655000 ;
      RECT 0.000000 240.465000 368.700000 240.615000 ;
      RECT 0.280000 240.235000 368.700000 240.465000 ;
      RECT 0.280000 240.085000 368.980000 240.235000 ;
      RECT 0.280000 240.045000 368.700000 240.085000 ;
      RECT 0.000000 239.895000 368.700000 240.045000 ;
      RECT 0.280000 239.665000 368.700000 239.895000 ;
      RECT 0.280000 239.515000 368.980000 239.665000 ;
      RECT 0.280000 239.475000 368.700000 239.515000 ;
      RECT 0.000000 239.325000 368.700000 239.475000 ;
      RECT 0.280000 239.095000 368.700000 239.325000 ;
      RECT 0.280000 238.945000 368.980000 239.095000 ;
      RECT 0.280000 238.905000 368.700000 238.945000 ;
      RECT 0.000000 238.755000 368.700000 238.905000 ;
      RECT 0.280000 238.525000 368.700000 238.755000 ;
      RECT 0.280000 238.375000 368.980000 238.525000 ;
      RECT 0.280000 238.335000 368.700000 238.375000 ;
      RECT 0.000000 238.185000 368.700000 238.335000 ;
      RECT 0.280000 237.955000 368.700000 238.185000 ;
      RECT 0.280000 237.805000 368.980000 237.955000 ;
      RECT 0.280000 237.765000 368.700000 237.805000 ;
      RECT 0.000000 237.615000 368.700000 237.765000 ;
      RECT 0.280000 237.385000 368.700000 237.615000 ;
      RECT 0.280000 237.235000 368.980000 237.385000 ;
      RECT 0.280000 237.195000 368.700000 237.235000 ;
      RECT 0.000000 237.045000 368.700000 237.195000 ;
      RECT 0.280000 236.815000 368.700000 237.045000 ;
      RECT 0.280000 236.665000 368.980000 236.815000 ;
      RECT 0.280000 236.625000 368.700000 236.665000 ;
      RECT 0.000000 236.475000 368.700000 236.625000 ;
      RECT 0.280000 236.245000 368.700000 236.475000 ;
      RECT 0.280000 236.095000 368.980000 236.245000 ;
      RECT 0.280000 236.055000 368.700000 236.095000 ;
      RECT 0.000000 235.905000 368.700000 236.055000 ;
      RECT 0.280000 235.675000 368.700000 235.905000 ;
      RECT 0.280000 235.525000 368.980000 235.675000 ;
      RECT 0.280000 235.485000 368.700000 235.525000 ;
      RECT 0.000000 235.335000 368.700000 235.485000 ;
      RECT 0.280000 235.105000 368.700000 235.335000 ;
      RECT 0.280000 234.955000 368.980000 235.105000 ;
      RECT 0.280000 234.915000 368.700000 234.955000 ;
      RECT 0.000000 234.765000 368.700000 234.915000 ;
      RECT 0.280000 234.535000 368.700000 234.765000 ;
      RECT 0.280000 234.385000 368.980000 234.535000 ;
      RECT 0.280000 234.345000 368.700000 234.385000 ;
      RECT 0.000000 234.195000 368.700000 234.345000 ;
      RECT 0.280000 233.965000 368.700000 234.195000 ;
      RECT 0.280000 233.815000 368.980000 233.965000 ;
      RECT 0.280000 233.775000 368.700000 233.815000 ;
      RECT 0.000000 233.625000 368.700000 233.775000 ;
      RECT 0.280000 233.395000 368.700000 233.625000 ;
      RECT 0.280000 233.245000 368.980000 233.395000 ;
      RECT 0.280000 233.205000 368.700000 233.245000 ;
      RECT 0.000000 233.055000 368.700000 233.205000 ;
      RECT 0.280000 232.825000 368.700000 233.055000 ;
      RECT 0.280000 232.675000 368.980000 232.825000 ;
      RECT 0.280000 232.635000 368.700000 232.675000 ;
      RECT 0.000000 232.485000 368.700000 232.635000 ;
      RECT 0.280000 232.255000 368.700000 232.485000 ;
      RECT 0.280000 232.105000 368.980000 232.255000 ;
      RECT 0.280000 232.065000 368.700000 232.105000 ;
      RECT 0.000000 231.915000 368.700000 232.065000 ;
      RECT 0.280000 231.685000 368.700000 231.915000 ;
      RECT 0.280000 231.535000 368.980000 231.685000 ;
      RECT 0.280000 231.495000 368.700000 231.535000 ;
      RECT 0.000000 231.345000 368.700000 231.495000 ;
      RECT 0.280000 231.115000 368.700000 231.345000 ;
      RECT 0.280000 230.965000 368.980000 231.115000 ;
      RECT 0.280000 230.925000 368.700000 230.965000 ;
      RECT 0.000000 230.775000 368.700000 230.925000 ;
      RECT 0.280000 230.545000 368.700000 230.775000 ;
      RECT 0.280000 230.395000 368.980000 230.545000 ;
      RECT 0.280000 230.355000 368.700000 230.395000 ;
      RECT 0.000000 230.205000 368.700000 230.355000 ;
      RECT 0.280000 229.975000 368.700000 230.205000 ;
      RECT 0.280000 229.825000 368.980000 229.975000 ;
      RECT 0.280000 229.785000 368.700000 229.825000 ;
      RECT 0.000000 229.635000 368.700000 229.785000 ;
      RECT 0.280000 229.405000 368.700000 229.635000 ;
      RECT 0.280000 229.255000 368.980000 229.405000 ;
      RECT 0.280000 229.215000 368.700000 229.255000 ;
      RECT 0.000000 229.065000 368.700000 229.215000 ;
      RECT 0.280000 228.835000 368.700000 229.065000 ;
      RECT 0.280000 228.685000 368.980000 228.835000 ;
      RECT 0.280000 228.645000 368.700000 228.685000 ;
      RECT 0.000000 228.495000 368.700000 228.645000 ;
      RECT 0.280000 228.265000 368.700000 228.495000 ;
      RECT 0.280000 228.115000 368.980000 228.265000 ;
      RECT 0.280000 228.075000 368.700000 228.115000 ;
      RECT 0.000000 227.925000 368.700000 228.075000 ;
      RECT 0.280000 227.695000 368.700000 227.925000 ;
      RECT 0.280000 227.545000 368.980000 227.695000 ;
      RECT 0.280000 227.505000 368.700000 227.545000 ;
      RECT 0.000000 227.355000 368.700000 227.505000 ;
      RECT 0.280000 227.125000 368.700000 227.355000 ;
      RECT 0.280000 226.975000 368.980000 227.125000 ;
      RECT 0.280000 226.935000 368.700000 226.975000 ;
      RECT 0.000000 226.785000 368.700000 226.935000 ;
      RECT 0.280000 226.555000 368.700000 226.785000 ;
      RECT 0.280000 226.405000 368.980000 226.555000 ;
      RECT 0.280000 226.365000 368.700000 226.405000 ;
      RECT 0.000000 226.215000 368.700000 226.365000 ;
      RECT 0.280000 225.985000 368.700000 226.215000 ;
      RECT 0.280000 225.835000 368.980000 225.985000 ;
      RECT 0.280000 225.795000 368.700000 225.835000 ;
      RECT 0.000000 225.645000 368.700000 225.795000 ;
      RECT 0.280000 225.415000 368.700000 225.645000 ;
      RECT 0.280000 225.265000 368.980000 225.415000 ;
      RECT 0.280000 225.225000 368.700000 225.265000 ;
      RECT 0.000000 225.075000 368.700000 225.225000 ;
      RECT 0.280000 224.845000 368.700000 225.075000 ;
      RECT 0.280000 224.695000 368.980000 224.845000 ;
      RECT 0.280000 224.655000 368.700000 224.695000 ;
      RECT 0.000000 224.505000 368.700000 224.655000 ;
      RECT 0.280000 224.275000 368.700000 224.505000 ;
      RECT 0.280000 224.125000 368.980000 224.275000 ;
      RECT 0.280000 224.085000 368.700000 224.125000 ;
      RECT 0.000000 223.935000 368.700000 224.085000 ;
      RECT 0.280000 223.705000 368.700000 223.935000 ;
      RECT 0.280000 223.555000 368.980000 223.705000 ;
      RECT 0.280000 223.515000 368.700000 223.555000 ;
      RECT 0.000000 223.365000 368.700000 223.515000 ;
      RECT 0.280000 223.135000 368.700000 223.365000 ;
      RECT 0.280000 222.985000 368.980000 223.135000 ;
      RECT 0.280000 222.945000 368.700000 222.985000 ;
      RECT 0.000000 222.795000 368.700000 222.945000 ;
      RECT 0.280000 222.565000 368.700000 222.795000 ;
      RECT 0.280000 222.415000 368.980000 222.565000 ;
      RECT 0.280000 222.375000 368.700000 222.415000 ;
      RECT 0.000000 222.225000 368.700000 222.375000 ;
      RECT 0.280000 221.995000 368.700000 222.225000 ;
      RECT 0.280000 221.845000 368.980000 221.995000 ;
      RECT 0.280000 221.805000 368.700000 221.845000 ;
      RECT 0.000000 221.655000 368.700000 221.805000 ;
      RECT 0.280000 221.425000 368.700000 221.655000 ;
      RECT 0.280000 221.275000 368.980000 221.425000 ;
      RECT 0.280000 221.235000 368.700000 221.275000 ;
      RECT 0.000000 221.085000 368.700000 221.235000 ;
      RECT 0.280000 220.855000 368.700000 221.085000 ;
      RECT 0.280000 220.705000 368.980000 220.855000 ;
      RECT 0.280000 220.665000 368.700000 220.705000 ;
      RECT 0.000000 220.515000 368.700000 220.665000 ;
      RECT 0.280000 220.285000 368.700000 220.515000 ;
      RECT 0.280000 220.135000 368.980000 220.285000 ;
      RECT 0.280000 220.095000 368.700000 220.135000 ;
      RECT 0.000000 219.945000 368.700000 220.095000 ;
      RECT 0.280000 219.715000 368.700000 219.945000 ;
      RECT 0.280000 219.565000 368.980000 219.715000 ;
      RECT 0.280000 219.525000 368.700000 219.565000 ;
      RECT 0.000000 219.375000 368.700000 219.525000 ;
      RECT 0.280000 219.145000 368.700000 219.375000 ;
      RECT 0.280000 218.995000 368.980000 219.145000 ;
      RECT 0.280000 218.955000 368.700000 218.995000 ;
      RECT 0.000000 218.805000 368.700000 218.955000 ;
      RECT 0.280000 218.575000 368.700000 218.805000 ;
      RECT 0.280000 218.425000 368.980000 218.575000 ;
      RECT 0.280000 218.385000 368.700000 218.425000 ;
      RECT 0.000000 218.235000 368.700000 218.385000 ;
      RECT 0.280000 218.005000 368.700000 218.235000 ;
      RECT 0.280000 217.855000 368.980000 218.005000 ;
      RECT 0.280000 217.815000 368.700000 217.855000 ;
      RECT 0.000000 217.665000 368.700000 217.815000 ;
      RECT 0.280000 217.435000 368.700000 217.665000 ;
      RECT 0.280000 217.285000 368.980000 217.435000 ;
      RECT 0.280000 217.245000 368.700000 217.285000 ;
      RECT 0.000000 217.095000 368.700000 217.245000 ;
      RECT 0.280000 216.865000 368.700000 217.095000 ;
      RECT 0.280000 216.715000 368.980000 216.865000 ;
      RECT 0.280000 216.675000 368.700000 216.715000 ;
      RECT 0.000000 216.525000 368.700000 216.675000 ;
      RECT 0.280000 216.295000 368.700000 216.525000 ;
      RECT 0.280000 216.145000 368.980000 216.295000 ;
      RECT 0.280000 216.105000 368.700000 216.145000 ;
      RECT 0.000000 215.955000 368.700000 216.105000 ;
      RECT 0.280000 215.725000 368.700000 215.955000 ;
      RECT 0.280000 215.575000 368.980000 215.725000 ;
      RECT 0.280000 215.535000 368.700000 215.575000 ;
      RECT 0.000000 215.385000 368.700000 215.535000 ;
      RECT 0.280000 215.155000 368.700000 215.385000 ;
      RECT 0.280000 215.005000 368.980000 215.155000 ;
      RECT 0.280000 214.965000 368.700000 215.005000 ;
      RECT 0.000000 214.815000 368.700000 214.965000 ;
      RECT 0.280000 214.585000 368.700000 214.815000 ;
      RECT 0.280000 214.435000 368.980000 214.585000 ;
      RECT 0.280000 214.395000 368.700000 214.435000 ;
      RECT 0.000000 214.245000 368.700000 214.395000 ;
      RECT 0.280000 214.015000 368.700000 214.245000 ;
      RECT 0.280000 213.865000 368.980000 214.015000 ;
      RECT 0.280000 213.825000 368.700000 213.865000 ;
      RECT 0.000000 213.675000 368.700000 213.825000 ;
      RECT 0.280000 213.445000 368.700000 213.675000 ;
      RECT 0.280000 213.295000 368.980000 213.445000 ;
      RECT 0.280000 213.255000 368.700000 213.295000 ;
      RECT 0.000000 213.105000 368.700000 213.255000 ;
      RECT 0.280000 212.875000 368.700000 213.105000 ;
      RECT 0.280000 212.725000 368.980000 212.875000 ;
      RECT 0.280000 212.685000 368.700000 212.725000 ;
      RECT 0.000000 212.535000 368.700000 212.685000 ;
      RECT 0.280000 212.305000 368.700000 212.535000 ;
      RECT 0.280000 212.155000 368.980000 212.305000 ;
      RECT 0.280000 212.115000 368.700000 212.155000 ;
      RECT 0.000000 211.965000 368.700000 212.115000 ;
      RECT 0.280000 211.735000 368.700000 211.965000 ;
      RECT 0.280000 211.585000 368.980000 211.735000 ;
      RECT 0.280000 211.545000 368.700000 211.585000 ;
      RECT 0.000000 211.395000 368.700000 211.545000 ;
      RECT 0.280000 211.165000 368.700000 211.395000 ;
      RECT 0.280000 211.015000 368.980000 211.165000 ;
      RECT 0.280000 210.975000 368.700000 211.015000 ;
      RECT 0.000000 210.825000 368.700000 210.975000 ;
      RECT 0.280000 210.595000 368.700000 210.825000 ;
      RECT 0.280000 210.445000 368.980000 210.595000 ;
      RECT 0.280000 210.405000 368.700000 210.445000 ;
      RECT 0.000000 210.255000 368.700000 210.405000 ;
      RECT 0.280000 210.025000 368.700000 210.255000 ;
      RECT 0.280000 209.875000 368.980000 210.025000 ;
      RECT 0.280000 209.835000 368.700000 209.875000 ;
      RECT 0.000000 209.685000 368.700000 209.835000 ;
      RECT 0.280000 209.455000 368.700000 209.685000 ;
      RECT 0.280000 209.305000 368.980000 209.455000 ;
      RECT 0.280000 209.265000 368.700000 209.305000 ;
      RECT 0.000000 209.115000 368.700000 209.265000 ;
      RECT 0.280000 208.885000 368.700000 209.115000 ;
      RECT 0.280000 208.735000 368.980000 208.885000 ;
      RECT 0.280000 208.695000 368.700000 208.735000 ;
      RECT 0.000000 208.545000 368.700000 208.695000 ;
      RECT 0.280000 208.315000 368.700000 208.545000 ;
      RECT 0.280000 208.165000 368.980000 208.315000 ;
      RECT 0.280000 208.125000 368.700000 208.165000 ;
      RECT 0.000000 207.975000 368.700000 208.125000 ;
      RECT 0.280000 207.745000 368.700000 207.975000 ;
      RECT 0.280000 207.595000 368.980000 207.745000 ;
      RECT 0.280000 207.555000 368.700000 207.595000 ;
      RECT 0.000000 207.405000 368.700000 207.555000 ;
      RECT 0.280000 207.175000 368.700000 207.405000 ;
      RECT 0.280000 207.025000 368.980000 207.175000 ;
      RECT 0.280000 206.985000 368.700000 207.025000 ;
      RECT 0.000000 206.835000 368.700000 206.985000 ;
      RECT 0.280000 206.605000 368.700000 206.835000 ;
      RECT 0.280000 206.455000 368.980000 206.605000 ;
      RECT 0.280000 206.415000 368.700000 206.455000 ;
      RECT 0.000000 206.265000 368.700000 206.415000 ;
      RECT 0.280000 206.035000 368.700000 206.265000 ;
      RECT 0.280000 205.885000 368.980000 206.035000 ;
      RECT 0.280000 205.845000 368.700000 205.885000 ;
      RECT 0.000000 205.695000 368.700000 205.845000 ;
      RECT 0.280000 205.465000 368.700000 205.695000 ;
      RECT 0.280000 205.315000 368.980000 205.465000 ;
      RECT 0.280000 205.275000 368.700000 205.315000 ;
      RECT 0.000000 205.125000 368.700000 205.275000 ;
      RECT 0.280000 204.895000 368.700000 205.125000 ;
      RECT 0.280000 204.745000 368.980000 204.895000 ;
      RECT 0.280000 204.705000 368.700000 204.745000 ;
      RECT 0.000000 204.555000 368.700000 204.705000 ;
      RECT 0.280000 204.325000 368.700000 204.555000 ;
      RECT 0.280000 204.175000 368.980000 204.325000 ;
      RECT 0.280000 204.135000 368.700000 204.175000 ;
      RECT 0.000000 203.985000 368.700000 204.135000 ;
      RECT 0.280000 203.755000 368.700000 203.985000 ;
      RECT 0.280000 203.605000 368.980000 203.755000 ;
      RECT 0.280000 203.565000 368.700000 203.605000 ;
      RECT 0.000000 203.415000 368.700000 203.565000 ;
      RECT 0.280000 203.185000 368.700000 203.415000 ;
      RECT 0.280000 203.035000 368.980000 203.185000 ;
      RECT 0.280000 202.995000 368.700000 203.035000 ;
      RECT 0.000000 202.845000 368.700000 202.995000 ;
      RECT 0.280000 202.615000 368.700000 202.845000 ;
      RECT 0.280000 202.465000 368.980000 202.615000 ;
      RECT 0.280000 202.425000 368.700000 202.465000 ;
      RECT 0.000000 202.275000 368.700000 202.425000 ;
      RECT 0.280000 202.045000 368.700000 202.275000 ;
      RECT 0.280000 201.895000 368.980000 202.045000 ;
      RECT 0.280000 201.855000 368.700000 201.895000 ;
      RECT 0.000000 201.705000 368.700000 201.855000 ;
      RECT 0.280000 201.475000 368.700000 201.705000 ;
      RECT 0.280000 201.325000 368.980000 201.475000 ;
      RECT 0.280000 201.285000 368.700000 201.325000 ;
      RECT 0.000000 201.135000 368.700000 201.285000 ;
      RECT 0.280000 200.905000 368.700000 201.135000 ;
      RECT 0.280000 200.755000 368.980000 200.905000 ;
      RECT 0.280000 200.715000 368.700000 200.755000 ;
      RECT 0.000000 200.565000 368.700000 200.715000 ;
      RECT 0.280000 200.335000 368.700000 200.565000 ;
      RECT 0.280000 200.185000 368.980000 200.335000 ;
      RECT 0.280000 200.145000 368.700000 200.185000 ;
      RECT 0.000000 199.995000 368.700000 200.145000 ;
      RECT 0.280000 199.765000 368.700000 199.995000 ;
      RECT 0.280000 199.615000 368.980000 199.765000 ;
      RECT 0.280000 199.575000 368.700000 199.615000 ;
      RECT 0.000000 199.425000 368.700000 199.575000 ;
      RECT 0.280000 199.195000 368.700000 199.425000 ;
      RECT 0.280000 199.045000 368.980000 199.195000 ;
      RECT 0.280000 199.005000 368.700000 199.045000 ;
      RECT 0.000000 198.855000 368.700000 199.005000 ;
      RECT 0.280000 198.625000 368.700000 198.855000 ;
      RECT 0.280000 198.475000 368.980000 198.625000 ;
      RECT 0.280000 198.435000 368.700000 198.475000 ;
      RECT 0.000000 198.285000 368.700000 198.435000 ;
      RECT 0.280000 198.055000 368.700000 198.285000 ;
      RECT 0.280000 197.905000 368.980000 198.055000 ;
      RECT 0.280000 197.865000 368.700000 197.905000 ;
      RECT 0.000000 197.715000 368.700000 197.865000 ;
      RECT 0.280000 197.485000 368.700000 197.715000 ;
      RECT 0.280000 197.335000 368.980000 197.485000 ;
      RECT 0.280000 197.295000 368.700000 197.335000 ;
      RECT 0.000000 197.145000 368.700000 197.295000 ;
      RECT 0.280000 196.915000 368.700000 197.145000 ;
      RECT 0.280000 196.765000 368.980000 196.915000 ;
      RECT 0.280000 196.725000 368.700000 196.765000 ;
      RECT 0.000000 196.575000 368.700000 196.725000 ;
      RECT 0.280000 196.345000 368.700000 196.575000 ;
      RECT 0.280000 196.195000 368.980000 196.345000 ;
      RECT 0.280000 196.155000 368.700000 196.195000 ;
      RECT 0.000000 196.005000 368.700000 196.155000 ;
      RECT 0.280000 195.775000 368.700000 196.005000 ;
      RECT 0.280000 195.625000 368.980000 195.775000 ;
      RECT 0.280000 195.585000 368.700000 195.625000 ;
      RECT 0.000000 195.435000 368.700000 195.585000 ;
      RECT 0.280000 195.205000 368.700000 195.435000 ;
      RECT 0.280000 195.055000 368.980000 195.205000 ;
      RECT 0.280000 195.015000 368.700000 195.055000 ;
      RECT 0.000000 194.865000 368.700000 195.015000 ;
      RECT 0.280000 194.635000 368.700000 194.865000 ;
      RECT 0.280000 194.485000 368.980000 194.635000 ;
      RECT 0.280000 194.445000 368.700000 194.485000 ;
      RECT 0.000000 194.295000 368.700000 194.445000 ;
      RECT 0.280000 194.065000 368.700000 194.295000 ;
      RECT 0.280000 193.915000 368.980000 194.065000 ;
      RECT 0.280000 193.875000 368.700000 193.915000 ;
      RECT 0.000000 193.725000 368.700000 193.875000 ;
      RECT 0.280000 193.495000 368.700000 193.725000 ;
      RECT 0.280000 193.345000 368.980000 193.495000 ;
      RECT 0.280000 193.305000 368.700000 193.345000 ;
      RECT 0.000000 193.155000 368.700000 193.305000 ;
      RECT 0.280000 192.925000 368.700000 193.155000 ;
      RECT 0.280000 192.775000 368.980000 192.925000 ;
      RECT 0.280000 192.735000 368.700000 192.775000 ;
      RECT 0.000000 192.585000 368.700000 192.735000 ;
      RECT 0.280000 192.355000 368.700000 192.585000 ;
      RECT 0.280000 192.205000 368.980000 192.355000 ;
      RECT 0.280000 192.165000 368.700000 192.205000 ;
      RECT 0.000000 192.015000 368.700000 192.165000 ;
      RECT 0.280000 191.785000 368.700000 192.015000 ;
      RECT 0.280000 191.635000 368.980000 191.785000 ;
      RECT 0.280000 191.595000 368.700000 191.635000 ;
      RECT 0.000000 191.445000 368.700000 191.595000 ;
      RECT 0.280000 191.215000 368.700000 191.445000 ;
      RECT 0.280000 191.065000 368.980000 191.215000 ;
      RECT 0.280000 191.025000 368.700000 191.065000 ;
      RECT 0.000000 190.875000 368.700000 191.025000 ;
      RECT 0.280000 190.645000 368.700000 190.875000 ;
      RECT 0.280000 190.495000 368.980000 190.645000 ;
      RECT 0.280000 190.455000 368.700000 190.495000 ;
      RECT 0.000000 190.305000 368.700000 190.455000 ;
      RECT 0.280000 190.075000 368.700000 190.305000 ;
      RECT 0.280000 189.925000 368.980000 190.075000 ;
      RECT 0.280000 189.885000 368.700000 189.925000 ;
      RECT 0.000000 189.735000 368.700000 189.885000 ;
      RECT 0.280000 189.505000 368.700000 189.735000 ;
      RECT 0.280000 189.355000 368.980000 189.505000 ;
      RECT 0.280000 189.315000 368.700000 189.355000 ;
      RECT 0.000000 189.165000 368.700000 189.315000 ;
      RECT 0.280000 188.935000 368.700000 189.165000 ;
      RECT 0.280000 188.785000 368.980000 188.935000 ;
      RECT 0.280000 188.745000 368.700000 188.785000 ;
      RECT 0.000000 188.595000 368.700000 188.745000 ;
      RECT 0.280000 188.365000 368.700000 188.595000 ;
      RECT 0.280000 188.215000 368.980000 188.365000 ;
      RECT 0.280000 188.175000 368.700000 188.215000 ;
      RECT 0.000000 188.025000 368.700000 188.175000 ;
      RECT 0.280000 187.795000 368.700000 188.025000 ;
      RECT 0.280000 187.645000 368.980000 187.795000 ;
      RECT 0.280000 187.605000 368.700000 187.645000 ;
      RECT 0.000000 187.455000 368.700000 187.605000 ;
      RECT 0.280000 187.225000 368.700000 187.455000 ;
      RECT 0.280000 187.075000 368.980000 187.225000 ;
      RECT 0.280000 187.035000 368.700000 187.075000 ;
      RECT 0.000000 186.885000 368.700000 187.035000 ;
      RECT 0.280000 186.655000 368.700000 186.885000 ;
      RECT 0.280000 186.505000 368.980000 186.655000 ;
      RECT 0.280000 186.465000 368.700000 186.505000 ;
      RECT 0.000000 186.315000 368.700000 186.465000 ;
      RECT 0.280000 186.085000 368.700000 186.315000 ;
      RECT 0.280000 185.935000 368.980000 186.085000 ;
      RECT 0.280000 185.895000 368.700000 185.935000 ;
      RECT 0.000000 185.745000 368.700000 185.895000 ;
      RECT 0.280000 185.515000 368.700000 185.745000 ;
      RECT 0.280000 185.365000 368.980000 185.515000 ;
      RECT 0.280000 185.325000 368.700000 185.365000 ;
      RECT 0.000000 185.175000 368.700000 185.325000 ;
      RECT 0.280000 184.945000 368.700000 185.175000 ;
      RECT 0.280000 184.795000 368.980000 184.945000 ;
      RECT 0.280000 184.755000 368.700000 184.795000 ;
      RECT 0.000000 184.605000 368.700000 184.755000 ;
      RECT 0.280000 184.375000 368.700000 184.605000 ;
      RECT 0.280000 184.225000 368.980000 184.375000 ;
      RECT 0.280000 184.185000 368.700000 184.225000 ;
      RECT 0.000000 184.035000 368.700000 184.185000 ;
      RECT 0.280000 183.805000 368.700000 184.035000 ;
      RECT 0.280000 183.655000 368.980000 183.805000 ;
      RECT 0.280000 183.615000 368.700000 183.655000 ;
      RECT 0.000000 183.465000 368.700000 183.615000 ;
      RECT 0.280000 183.235000 368.700000 183.465000 ;
      RECT 0.280000 183.085000 368.980000 183.235000 ;
      RECT 0.280000 183.045000 368.700000 183.085000 ;
      RECT 0.000000 182.895000 368.700000 183.045000 ;
      RECT 0.280000 182.665000 368.700000 182.895000 ;
      RECT 0.280000 182.515000 368.980000 182.665000 ;
      RECT 0.280000 182.475000 368.700000 182.515000 ;
      RECT 0.000000 182.325000 368.700000 182.475000 ;
      RECT 0.280000 182.095000 368.700000 182.325000 ;
      RECT 0.280000 181.945000 368.980000 182.095000 ;
      RECT 0.280000 181.905000 368.700000 181.945000 ;
      RECT 0.000000 181.755000 368.700000 181.905000 ;
      RECT 0.280000 181.525000 368.700000 181.755000 ;
      RECT 0.280000 181.375000 368.980000 181.525000 ;
      RECT 0.280000 181.335000 368.700000 181.375000 ;
      RECT 0.000000 181.185000 368.700000 181.335000 ;
      RECT 0.280000 180.955000 368.700000 181.185000 ;
      RECT 0.280000 180.805000 368.980000 180.955000 ;
      RECT 0.280000 180.765000 368.700000 180.805000 ;
      RECT 0.000000 180.615000 368.700000 180.765000 ;
      RECT 0.280000 180.385000 368.700000 180.615000 ;
      RECT 0.280000 180.235000 368.980000 180.385000 ;
      RECT 0.280000 180.195000 368.700000 180.235000 ;
      RECT 0.000000 180.045000 368.700000 180.195000 ;
      RECT 0.280000 179.815000 368.700000 180.045000 ;
      RECT 0.280000 179.665000 368.980000 179.815000 ;
      RECT 0.280000 179.625000 368.700000 179.665000 ;
      RECT 0.000000 179.475000 368.700000 179.625000 ;
      RECT 0.280000 179.245000 368.700000 179.475000 ;
      RECT 0.280000 179.095000 368.980000 179.245000 ;
      RECT 0.280000 179.055000 368.700000 179.095000 ;
      RECT 0.000000 178.905000 368.700000 179.055000 ;
      RECT 0.280000 178.675000 368.700000 178.905000 ;
      RECT 0.280000 178.525000 368.980000 178.675000 ;
      RECT 0.280000 178.485000 368.700000 178.525000 ;
      RECT 0.000000 178.335000 368.700000 178.485000 ;
      RECT 0.280000 178.105000 368.700000 178.335000 ;
      RECT 0.280000 177.955000 368.980000 178.105000 ;
      RECT 0.280000 177.915000 368.700000 177.955000 ;
      RECT 0.000000 177.765000 368.700000 177.915000 ;
      RECT 0.280000 177.535000 368.700000 177.765000 ;
      RECT 0.280000 177.385000 368.980000 177.535000 ;
      RECT 0.280000 177.345000 368.700000 177.385000 ;
      RECT 0.000000 177.195000 368.700000 177.345000 ;
      RECT 0.280000 176.965000 368.700000 177.195000 ;
      RECT 0.280000 176.815000 368.980000 176.965000 ;
      RECT 0.280000 176.775000 368.700000 176.815000 ;
      RECT 0.000000 176.625000 368.700000 176.775000 ;
      RECT 0.280000 176.395000 368.700000 176.625000 ;
      RECT 0.280000 176.245000 368.980000 176.395000 ;
      RECT 0.280000 176.205000 368.700000 176.245000 ;
      RECT 0.000000 176.055000 368.700000 176.205000 ;
      RECT 0.280000 175.825000 368.700000 176.055000 ;
      RECT 0.280000 175.675000 368.980000 175.825000 ;
      RECT 0.280000 175.635000 368.700000 175.675000 ;
      RECT 0.000000 175.485000 368.700000 175.635000 ;
      RECT 0.280000 175.255000 368.700000 175.485000 ;
      RECT 0.280000 175.105000 368.980000 175.255000 ;
      RECT 0.280000 175.065000 368.700000 175.105000 ;
      RECT 0.000000 174.915000 368.700000 175.065000 ;
      RECT 0.280000 174.685000 368.700000 174.915000 ;
      RECT 0.280000 174.535000 368.980000 174.685000 ;
      RECT 0.280000 174.495000 368.700000 174.535000 ;
      RECT 0.000000 174.345000 368.700000 174.495000 ;
      RECT 0.280000 174.115000 368.700000 174.345000 ;
      RECT 0.280000 173.965000 368.980000 174.115000 ;
      RECT 0.280000 173.925000 368.700000 173.965000 ;
      RECT 0.000000 173.775000 368.700000 173.925000 ;
      RECT 0.280000 173.545000 368.700000 173.775000 ;
      RECT 0.280000 173.355000 368.980000 173.545000 ;
      RECT 0.000000 173.205000 368.980000 173.355000 ;
      RECT 0.280000 172.785000 368.980000 173.205000 ;
      RECT 0.000000 172.635000 368.980000 172.785000 ;
      RECT 0.280000 172.215000 368.980000 172.635000 ;
      RECT 0.000000 172.065000 368.980000 172.215000 ;
      RECT 0.280000 171.645000 368.980000 172.065000 ;
      RECT 0.000000 171.495000 368.980000 171.645000 ;
      RECT 0.280000 171.075000 368.980000 171.495000 ;
      RECT 0.000000 170.925000 368.980000 171.075000 ;
      RECT 0.280000 170.505000 368.980000 170.925000 ;
      RECT 0.000000 170.355000 368.980000 170.505000 ;
      RECT 0.280000 169.935000 368.980000 170.355000 ;
      RECT 0.000000 169.785000 368.980000 169.935000 ;
      RECT 0.280000 169.365000 368.980000 169.785000 ;
      RECT 0.000000 169.215000 368.980000 169.365000 ;
      RECT 0.280000 168.795000 368.980000 169.215000 ;
      RECT 0.000000 168.645000 368.980000 168.795000 ;
      RECT 0.280000 168.225000 368.980000 168.645000 ;
      RECT 0.000000 168.075000 368.980000 168.225000 ;
      RECT 0.280000 167.655000 368.980000 168.075000 ;
      RECT 0.000000 167.505000 368.980000 167.655000 ;
      RECT 0.280000 167.085000 368.980000 167.505000 ;
      RECT 0.000000 166.935000 368.980000 167.085000 ;
      RECT 0.280000 166.515000 368.980000 166.935000 ;
      RECT 0.000000 166.365000 368.980000 166.515000 ;
      RECT 0.280000 165.945000 368.980000 166.365000 ;
      RECT 0.000000 165.795000 368.980000 165.945000 ;
      RECT 0.280000 165.375000 368.980000 165.795000 ;
      RECT 0.000000 165.225000 368.980000 165.375000 ;
      RECT 0.280000 164.805000 368.980000 165.225000 ;
      RECT 0.000000 164.655000 368.980000 164.805000 ;
      RECT 0.280000 164.235000 368.980000 164.655000 ;
      RECT 0.000000 164.085000 368.980000 164.235000 ;
      RECT 0.280000 163.665000 368.980000 164.085000 ;
      RECT 0.000000 163.515000 368.980000 163.665000 ;
      RECT 0.280000 163.095000 368.980000 163.515000 ;
      RECT 0.000000 162.945000 368.980000 163.095000 ;
      RECT 0.280000 162.525000 368.980000 162.945000 ;
      RECT 0.000000 162.375000 368.980000 162.525000 ;
      RECT 0.280000 161.955000 368.980000 162.375000 ;
      RECT 0.000000 161.805000 368.980000 161.955000 ;
      RECT 0.280000 161.385000 368.980000 161.805000 ;
      RECT 0.000000 161.235000 368.980000 161.385000 ;
      RECT 0.280000 160.815000 368.980000 161.235000 ;
      RECT 0.000000 160.665000 368.980000 160.815000 ;
      RECT 0.280000 160.245000 368.980000 160.665000 ;
      RECT 0.000000 160.095000 368.980000 160.245000 ;
      RECT 0.280000 159.675000 368.980000 160.095000 ;
      RECT 0.000000 159.525000 368.980000 159.675000 ;
      RECT 0.280000 159.105000 368.980000 159.525000 ;
      RECT 0.000000 158.955000 368.980000 159.105000 ;
      RECT 0.280000 158.535000 368.980000 158.955000 ;
      RECT 0.000000 158.385000 368.980000 158.535000 ;
      RECT 0.280000 157.965000 368.980000 158.385000 ;
      RECT 0.000000 157.815000 368.980000 157.965000 ;
      RECT 0.280000 157.395000 368.980000 157.815000 ;
      RECT 0.000000 157.245000 368.980000 157.395000 ;
      RECT 0.280000 156.825000 368.980000 157.245000 ;
      RECT 0.000000 156.675000 368.980000 156.825000 ;
      RECT 0.280000 156.255000 368.980000 156.675000 ;
      RECT 0.000000 156.105000 368.980000 156.255000 ;
      RECT 0.280000 155.685000 368.980000 156.105000 ;
      RECT 0.000000 155.535000 368.980000 155.685000 ;
      RECT 0.280000 155.115000 368.980000 155.535000 ;
      RECT 0.000000 154.965000 368.980000 155.115000 ;
      RECT 0.280000 154.545000 368.980000 154.965000 ;
      RECT 0.000000 154.395000 368.980000 154.545000 ;
      RECT 0.280000 153.975000 368.980000 154.395000 ;
      RECT 0.000000 153.825000 368.980000 153.975000 ;
      RECT 0.280000 153.405000 368.980000 153.825000 ;
      RECT 0.000000 153.255000 368.980000 153.405000 ;
      RECT 0.280000 152.835000 368.980000 153.255000 ;
      RECT 0.000000 152.685000 368.980000 152.835000 ;
      RECT 0.280000 152.265000 368.980000 152.685000 ;
      RECT 0.000000 152.115000 368.980000 152.265000 ;
      RECT 0.280000 151.695000 368.980000 152.115000 ;
      RECT 0.000000 151.545000 368.980000 151.695000 ;
      RECT 0.280000 151.125000 368.980000 151.545000 ;
      RECT 0.000000 150.975000 368.980000 151.125000 ;
      RECT 0.280000 150.555000 368.980000 150.975000 ;
      RECT 0.000000 150.405000 368.980000 150.555000 ;
      RECT 0.280000 149.985000 368.980000 150.405000 ;
      RECT 0.000000 149.835000 368.980000 149.985000 ;
      RECT 0.280000 149.415000 368.980000 149.835000 ;
      RECT 0.000000 149.265000 368.980000 149.415000 ;
      RECT 0.280000 148.845000 368.980000 149.265000 ;
      RECT 0.000000 148.695000 368.980000 148.845000 ;
      RECT 0.280000 148.275000 368.980000 148.695000 ;
      RECT 0.000000 148.125000 368.980000 148.275000 ;
      RECT 0.280000 147.705000 368.980000 148.125000 ;
      RECT 0.000000 147.555000 368.980000 147.705000 ;
      RECT 0.280000 147.135000 368.980000 147.555000 ;
      RECT 0.000000 146.985000 368.980000 147.135000 ;
      RECT 0.280000 146.565000 368.980000 146.985000 ;
      RECT 0.000000 146.415000 368.980000 146.565000 ;
      RECT 0.280000 145.995000 368.980000 146.415000 ;
      RECT 0.000000 145.845000 368.980000 145.995000 ;
      RECT 0.280000 145.425000 368.980000 145.845000 ;
      RECT 0.000000 145.275000 368.980000 145.425000 ;
      RECT 0.280000 144.855000 368.980000 145.275000 ;
      RECT 0.000000 144.705000 368.980000 144.855000 ;
      RECT 0.280000 144.285000 368.980000 144.705000 ;
      RECT 0.000000 0.280000 368.980000 144.285000 ;
      RECT 21.865000 0.000000 368.980000 0.280000 ;
      RECT 20.185000 0.000000 21.445000 0.280000 ;
      RECT 18.225000 0.000000 19.765000 0.280000 ;
      RECT 16.545000 0.000000 17.805000 0.280000 ;
      RECT 14.585000 0.000000 16.125000 0.280000 ;
      RECT 12.625000 0.000000 14.165000 0.280000 ;
      RECT 10.945000 0.000000 12.205000 0.280000 ;
      RECT 8.985000 0.000000 10.525000 0.280000 ;
      RECT 7.025000 0.000000 8.565000 0.280000 ;
      RECT 5.345000 0.000000 6.605000 0.280000 ;
      RECT 0.000000 0.000000 4.925000 0.280000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 368.980000 437.570000 ;
  END
END MLP_no_sram

END LIBRARY
