module SigmoidTable(
	input [15:0] x,
	output reg [7:0] y
);

always @(*) begin
	if(x[15:7]==9'h1FF || x[15:7]==9'h000)begin
		case(x[7:0])
			8'h00 : y = 8'h10;		// Float Value -> 0.5
			8'h01 : y = 8'h10;		// Float Value -> 0.5
			8'h02 : y = 8'h10;		// Float Value -> 0.5
			8'h03 : y = 8'h10;		// Float Value -> 0.5
			8'h04 : y = 8'h10;		// Float Value -> 0.5
			8'h05 : y = 8'h11;		// Float Value -> 0.53125
			8'h06 : y = 8'h11;		// Float Value -> 0.53125
			8'h07 : y = 8'h11;		// Float Value -> 0.53125
			8'h08 : y = 8'h11;		// Float Value -> 0.53125
			8'h09 : y = 8'h12;		// Float Value -> 0.5625
			8'h0A : y = 8'h12;		// Float Value -> 0.5625
			8'h0B : y = 8'h12;		// Float Value -> 0.5625
			8'h0C : y = 8'h12;		// Float Value -> 0.5625
			8'h0D : y = 8'h13;		// Float Value -> 0.59375
			8'h0E : y = 8'h13;		// Float Value -> 0.59375
			8'h0F : y = 8'h13;		// Float Value -> 0.59375
			8'h10 : y = 8'h13;		// Float Value -> 0.59375
			8'h11 : y = 8'h14;		// Float Value -> 0.625
			8'h12 : y = 8'h14;		// Float Value -> 0.625
			8'h13 : y = 8'h14;		// Float Value -> 0.625
			8'h14 : y = 8'h14;		// Float Value -> 0.625
			8'h15 : y = 8'h15;		// Float Value -> 0.65625
			8'h16 : y = 8'h15;		// Float Value -> 0.65625
			8'h17 : y = 8'h15;		// Float Value -> 0.65625
			8'h18 : y = 8'h15;		// Float Value -> 0.65625
			8'h19 : y = 8'h15;		// Float Value -> 0.65625
			8'h1A : y = 8'h16;		// Float Value -> 0.6875
			8'h1B : y = 8'h16;		// Float Value -> 0.6875
			8'h1C : y = 8'h16;		// Float Value -> 0.6875
			8'h1D : y = 8'h16;		// Float Value -> 0.6875
			8'h1E : y = 8'h16;		// Float Value -> 0.6875
			8'h1F : y = 8'h17;		// Float Value -> 0.71875
			8'h20 : y = 8'h17;		// Float Value -> 0.71875
			8'h21 : y = 8'h17;		// Float Value -> 0.71875
			8'h22 : y = 8'h17;		// Float Value -> 0.71875
			8'h23 : y = 8'h17;		// Float Value -> 0.71875
			8'h24 : y = 8'h18;		// Float Value -> 0.75
			8'h25 : y = 8'h18;		// Float Value -> 0.75
			8'h26 : y = 8'h18;		// Float Value -> 0.75
			8'h27 : y = 8'h18;		// Float Value -> 0.75
			8'h28 : y = 8'h18;		// Float Value -> 0.75
			8'h29 : y = 8'h19;		// Float Value -> 0.78125
			8'h2A : y = 8'h19;		// Float Value -> 0.78125
			8'h2B : y = 8'h19;		// Float Value -> 0.78125
			8'h2C : y = 8'h19;		// Float Value -> 0.78125
			8'h2D : y = 8'h19;		// Float Value -> 0.78125
			8'h2E : y = 8'h19;		// Float Value -> 0.78125
			8'h2F : y = 8'h1A;		// Float Value -> 0.8125
			8'h30 : y = 8'h1A;		// Float Value -> 0.8125
			8'h31 : y = 8'h1A;		// Float Value -> 0.8125
			8'h32 : y = 8'h1A;		// Float Value -> 0.8125
			8'h33 : y = 8'h1A;		// Float Value -> 0.8125
			8'h34 : y = 8'h1A;		// Float Value -> 0.8125
			8'h35 : y = 8'h1A;		// Float Value -> 0.8125
			8'h36 : y = 8'h1B;		// Float Value -> 0.84375
			8'h37 : y = 8'h1B;		// Float Value -> 0.84375
			8'h38 : y = 8'h1B;		// Float Value -> 0.84375
			8'h39 : y = 8'h1B;		// Float Value -> 0.84375
			8'h3A : y = 8'h1B;		// Float Value -> 0.84375
			8'h3B : y = 8'h1B;		// Float Value -> 0.84375
			8'h3C : y = 8'h1B;		// Float Value -> 0.84375
			8'h3D : y = 8'h1B;		// Float Value -> 0.84375
			8'h3E : y = 8'h1B;		// Float Value -> 0.84375
			8'h3F : y = 8'h1C;		// Float Value -> 0.875
			8'h40 : y = 8'h1C;		// Float Value -> 0.875
			8'h41 : y = 8'h1C;		// Float Value -> 0.875
			8'h42 : y = 8'h1C;		// Float Value -> 0.875
			8'h43 : y = 8'h1C;		// Float Value -> 0.875
			8'h44 : y = 8'h1C;		// Float Value -> 0.875
			8'h45 : y = 8'h1C;		// Float Value -> 0.875
			8'h46 : y = 8'h1C;		// Float Value -> 0.875
			8'h47 : y = 8'h1C;		// Float Value -> 0.875
			8'h48 : y = 8'h1C;		// Float Value -> 0.875
			8'h49 : y = 8'h1D;		// Float Value -> 0.90625
			8'h4A : y = 8'h1D;		// Float Value -> 0.90625
			8'h4B : y = 8'h1D;		// Float Value -> 0.90625
			8'h4C : y = 8'h1D;		// Float Value -> 0.90625
			8'h4D : y = 8'h1D;		// Float Value -> 0.90625
			8'h4E : y = 8'h1D;		// Float Value -> 0.90625
			8'h4F : y = 8'h1D;		// Float Value -> 0.90625
			8'h50 : y = 8'h1D;		// Float Value -> 0.90625
			8'h51 : y = 8'h1D;		// Float Value -> 0.90625
			8'h52 : y = 8'h1D;		// Float Value -> 0.90625
			8'h53 : y = 8'h1D;		// Float Value -> 0.90625
			8'h54 : y = 8'h1D;		// Float Value -> 0.90625
			8'h55 : y = 8'h1D;		// Float Value -> 0.90625
			8'h56 : y = 8'h1D;		// Float Value -> 0.90625
			8'h57 : y = 8'h1E;		// Float Value -> 0.9375
			8'h58 : y = 8'h1E;		// Float Value -> 0.9375
			8'h59 : y = 8'h1E;		// Float Value -> 0.9375
			8'h5A : y = 8'h1E;		// Float Value -> 0.9375
			8'h5B : y = 8'h1E;		// Float Value -> 0.9375
			8'h5C : y = 8'h1E;		// Float Value -> 0.9375
			8'h5D : y = 8'h1E;		// Float Value -> 0.9375
			8'h5E : y = 8'h1E;		// Float Value -> 0.9375
			8'h5F : y = 8'h1E;		// Float Value -> 0.9375
			8'h60 : y = 8'h1E;		// Float Value -> 0.9375
			8'h61 : y = 8'h1E;		// Float Value -> 0.9375
			8'h62 : y = 8'h1E;		// Float Value -> 0.9375
			8'h63 : y = 8'h1E;		// Float Value -> 0.9375
			8'h64 : y = 8'h1E;		// Float Value -> 0.9375
			8'h65 : y = 8'h1E;		// Float Value -> 0.9375
			8'h66 : y = 8'h1E;		// Float Value -> 0.9375
			8'h67 : y = 8'h1E;		// Float Value -> 0.9375
			8'h68 : y = 8'h1E;		// Float Value -> 0.9375
			8'h69 : y = 8'h1E;		// Float Value -> 0.9375
			8'h6A : y = 8'h1E;		// Float Value -> 0.9375
			8'h6B : y = 8'h1E;		// Float Value -> 0.9375
			8'h6C : y = 8'h1E;		// Float Value -> 0.9375
			8'h6D : y = 8'h1E;		// Float Value -> 0.9375
			8'h6E : y = 8'h1F;		// Float Value -> 0.96875
			8'h6F : y = 8'h1F;		// Float Value -> 0.96875
			8'h70 : y = 8'h1F;		// Float Value -> 0.96875
			8'h71 : y = 8'h1F;		// Float Value -> 0.96875
			8'h72 : y = 8'h1F;		// Float Value -> 0.96875
			8'h73 : y = 8'h1F;		// Float Value -> 0.96875
			8'h74 : y = 8'h1F;		// Float Value -> 0.96875
			8'h75 : y = 8'h1F;		// Float Value -> 0.96875
			8'h76 : y = 8'h1F;		// Float Value -> 0.96875
			8'h77 : y = 8'h1F;		// Float Value -> 0.96875
			8'h78 : y = 8'h1F;		// Float Value -> 0.96875
			8'h79 : y = 8'h1F;		// Float Value -> 0.96875
			8'h7A : y = 8'h1F;		// Float Value -> 0.96875
			8'h7B : y = 8'h1F;		// Float Value -> 0.96875
			8'h7C : y = 8'h1F;		// Float Value -> 0.96875
			8'h7D : y = 8'h1F;		// Float Value -> 0.96875
			8'h7E : y = 8'h1F;		// Float Value -> 0.96875
			8'h7F : y = 8'h1F;		// Float Value -> 0.96875
			8'h80 : y = 8'h00;		// Float Value -> 0.0
			8'h81 : y = 8'h00;		// Float Value -> 0.0
			8'h82 : y = 8'h00;		// Float Value -> 0.0
			8'h83 : y = 8'h00;		// Float Value -> 0.0
			8'h84 : y = 8'h00;		// Float Value -> 0.0
			8'h85 : y = 8'h00;		// Float Value -> 0.0
			8'h86 : y = 8'h00;		// Float Value -> 0.0
			8'h87 : y = 8'h00;		// Float Value -> 0.0
			8'h88 : y = 8'h00;		// Float Value -> 0.0
			8'h89 : y = 8'h00;		// Float Value -> 0.0
			8'h8A : y = 8'h00;		// Float Value -> 0.0
			8'h8B : y = 8'h00;		// Float Value -> 0.0
			8'h8C : y = 8'h00;		// Float Value -> 0.0
			8'h8D : y = 8'h00;		// Float Value -> 0.0
			8'h8E : y = 8'h00;		// Float Value -> 0.0
			8'h8F : y = 8'h00;		// Float Value -> 0.0
			8'h90 : y = 8'h00;		// Float Value -> 0.0
			8'h91 : y = 8'h00;		// Float Value -> 0.0
			8'h92 : y = 8'h00;		// Float Value -> 0.0
			8'h93 : y = 8'h01;		// Float Value -> 0.03125
			8'h94 : y = 8'h01;		// Float Value -> 0.03125
			8'h95 : y = 8'h01;		// Float Value -> 0.03125
			8'h96 : y = 8'h01;		// Float Value -> 0.03125
			8'h97 : y = 8'h01;		// Float Value -> 0.03125
			8'h98 : y = 8'h01;		// Float Value -> 0.03125
			8'h99 : y = 8'h01;		// Float Value -> 0.03125
			8'h9A : y = 8'h01;		// Float Value -> 0.03125
			8'h9B : y = 8'h01;		// Float Value -> 0.03125
			8'h9C : y = 8'h01;		// Float Value -> 0.03125
			8'h9D : y = 8'h01;		// Float Value -> 0.03125
			8'h9E : y = 8'h01;		// Float Value -> 0.03125
			8'h9F : y = 8'h01;		// Float Value -> 0.03125
			8'hA0 : y = 8'h01;		// Float Value -> 0.03125
			8'hA1 : y = 8'h01;		// Float Value -> 0.03125
			8'hA2 : y = 8'h01;		// Float Value -> 0.03125
			8'hA3 : y = 8'h01;		// Float Value -> 0.03125
			8'hA4 : y = 8'h01;		// Float Value -> 0.03125
			8'hA5 : y = 8'h01;		// Float Value -> 0.03125
			8'hA6 : y = 8'h01;		// Float Value -> 0.03125
			8'hA7 : y = 8'h01;		// Float Value -> 0.03125
			8'hA8 : y = 8'h01;		// Float Value -> 0.03125
			8'hA9 : y = 8'h01;		// Float Value -> 0.03125
			8'hAA : y = 8'h02;		// Float Value -> 0.0625
			8'hAB : y = 8'h02;		// Float Value -> 0.0625
			8'hAC : y = 8'h02;		// Float Value -> 0.0625
			8'hAD : y = 8'h02;		// Float Value -> 0.0625
			8'hAE : y = 8'h02;		// Float Value -> 0.0625
			8'hAF : y = 8'h02;		// Float Value -> 0.0625
			8'hB0 : y = 8'h02;		// Float Value -> 0.0625
			8'hB1 : y = 8'h02;		// Float Value -> 0.0625
			8'hB2 : y = 8'h02;		// Float Value -> 0.0625
			8'hB3 : y = 8'h02;		// Float Value -> 0.0625
			8'hB4 : y = 8'h02;		// Float Value -> 0.0625
			8'hB5 : y = 8'h02;		// Float Value -> 0.0625
			8'hB6 : y = 8'h02;		// Float Value -> 0.0625
			8'hB7 : y = 8'h02;		// Float Value -> 0.0625
			8'hB8 : y = 8'h03;		// Float Value -> 0.09375
			8'hB9 : y = 8'h03;		// Float Value -> 0.09375
			8'hBA : y = 8'h03;		// Float Value -> 0.09375
			8'hBB : y = 8'h03;		// Float Value -> 0.09375
			8'hBC : y = 8'h03;		// Float Value -> 0.09375
			8'hBD : y = 8'h03;		// Float Value -> 0.09375
			8'hBE : y = 8'h03;		// Float Value -> 0.09375
			8'hBF : y = 8'h03;		// Float Value -> 0.09375
			8'hC0 : y = 8'h03;		// Float Value -> 0.09375
			8'hC1 : y = 8'h03;		// Float Value -> 0.09375
			8'hC2 : y = 8'h04;		// Float Value -> 0.125
			8'hC3 : y = 8'h04;		// Float Value -> 0.125
			8'hC4 : y = 8'h04;		// Float Value -> 0.125
			8'hC5 : y = 8'h04;		// Float Value -> 0.125
			8'hC6 : y = 8'h04;		// Float Value -> 0.125
			8'hC7 : y = 8'h04;		// Float Value -> 0.125
			8'hC8 : y = 8'h04;		// Float Value -> 0.125
			8'hC9 : y = 8'h04;		// Float Value -> 0.125
			8'hCA : y = 8'h04;		// Float Value -> 0.125
			8'hCB : y = 8'h05;		// Float Value -> 0.15625
			8'hCC : y = 8'h05;		// Float Value -> 0.15625
			8'hCD : y = 8'h05;		// Float Value -> 0.15625
			8'hCE : y = 8'h05;		// Float Value -> 0.15625
			8'hCF : y = 8'h05;		// Float Value -> 0.15625
			8'hD0 : y = 8'h05;		// Float Value -> 0.15625
			8'hD1 : y = 8'h05;		// Float Value -> 0.15625
			8'hD2 : y = 8'h06;		// Float Value -> 0.1875
			8'hD3 : y = 8'h06;		// Float Value -> 0.1875
			8'hD4 : y = 8'h06;		// Float Value -> 0.1875
			8'hD5 : y = 8'h06;		// Float Value -> 0.1875
			8'hD6 : y = 8'h06;		// Float Value -> 0.1875
			8'hD7 : y = 8'h06;		// Float Value -> 0.1875
			8'hD8 : y = 8'h07;		// Float Value -> 0.21875
			8'hD9 : y = 8'h07;		// Float Value -> 0.21875
			8'hDA : y = 8'h07;		// Float Value -> 0.21875
			8'hDB : y = 8'h07;		// Float Value -> 0.21875
			8'hDC : y = 8'h07;		// Float Value -> 0.21875
			8'hDD : y = 8'h08;		// Float Value -> 0.25
			8'hDE : y = 8'h08;		// Float Value -> 0.25
			8'hDF : y = 8'h08;		// Float Value -> 0.25
			8'hE0 : y = 8'h08;		// Float Value -> 0.25
			8'hE1 : y = 8'h08;		// Float Value -> 0.25
			8'hE2 : y = 8'h09;		// Float Value -> 0.28125
			8'hE3 : y = 8'h09;		// Float Value -> 0.28125
			8'hE4 : y = 8'h09;		// Float Value -> 0.28125
			8'hE5 : y = 8'h09;		// Float Value -> 0.28125
			8'hE6 : y = 8'h09;		// Float Value -> 0.28125
			8'hE7 : y = 8'h0A;		// Float Value -> 0.3125
			8'hE8 : y = 8'h0A;		// Float Value -> 0.3125
			8'hE9 : y = 8'h0A;		// Float Value -> 0.3125
			8'hEA : y = 8'h0A;		// Float Value -> 0.3125
			8'hEB : y = 8'h0A;		// Float Value -> 0.3125
			8'hEC : y = 8'h0B;		// Float Value -> 0.34375
			8'hED : y = 8'h0B;		// Float Value -> 0.34375
			8'hEE : y = 8'h0B;		// Float Value -> 0.34375
			8'hEF : y = 8'h0B;		// Float Value -> 0.34375
			8'hF0 : y = 8'h0C;		// Float Value -> 0.375
			8'hF1 : y = 8'h0C;		// Float Value -> 0.375
			8'hF2 : y = 8'h0C;		// Float Value -> 0.375
			8'hF3 : y = 8'h0C;		// Float Value -> 0.375
			8'hF4 : y = 8'h0D;		// Float Value -> 0.40625
			8'hF5 : y = 8'h0D;		// Float Value -> 0.40625
			8'hF6 : y = 8'h0D;		// Float Value -> 0.40625
			8'hF7 : y = 8'h0D;		// Float Value -> 0.40625
			8'hF8 : y = 8'h0E;		// Float Value -> 0.4375
			8'hF9 : y = 8'h0E;		// Float Value -> 0.4375
			8'hFA : y = 8'h0E;		// Float Value -> 0.4375
			8'hFB : y = 8'h0E;		// Float Value -> 0.4375
			8'hFC : y = 8'h0F;		// Float Value -> 0.46875
			8'hFD : y = 8'h0F;		// Float Value -> 0.46875
			8'hFE : y = 8'h0F;		// Float Value -> 0.46875
			8'hFF : y = 8'h0F;		// Float Value -> 0.46875
			default : y = 8'h00;
		endcase
	end
	else begin
		if(x[15])begin
			y = 8'h00;
		end	
		else begin 		
			y = 8'h20;
		end
	end
end
endmodule
